///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: tf_ROM.v
// File history:
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// <Description here>
//
// Targeted device: <Family::PolarFireSoC> <Die::MPFS250T_ES> <Package::FCVG484>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

//`timescale <time_units> / <precision>

module tf0_ROM (
    input                       clk,
    input      [5:0]            A,
    output reg [11:0]           Q
);
    
    always@(posedge clk) begin
        case(A)
            6'd0: Q <= 12'd1201;
            6'd1: Q <= 12'd1434;
            6'd2: Q <= 12'd2610;
            6'd3: Q <= 12'd2382;
            6'd4: Q <= 12'd505;
            6'd5: Q <= 12'd226;
            6'd6: Q <= 12'd1261;
            6'd7: Q <= 12'd2278;
            6'd8: Q <= 12'd455;
            6'd9: Q <= 12'd1555;
            6'd10: Q <= 12'd2092;
            6'd11: Q <= 12'd2973;
            6'd12: Q <= 12'd341;
            6'd13: Q <= 12'd324;
            6'd14: Q <= 12'd924;
            6'd15: Q <= 12'd660;
            6'd16: Q <= 12'd2622;
            6'd17: Q <= 12'd1681;
            6'd18: Q <= 12'd232;
            6'd19: Q <= 12'd2653;
            6'd20: Q <= 12'd3004;
            6'd21: Q <= 12'd316;
            6'd22: Q <= 12'd408;
            6'd23: Q <= 12'd1830;
            6'd24: Q <= 12'd1520;
            6'd25: Q <= 12'd878;
            6'd26: Q <= 12'd38;
            6'd27: Q <= 12'd1152;
            6'd28: Q <= 12'd1066;
            6'd29: Q <= 12'd2692;
            6'd30: Q <= 12'd526;
            6'd31: Q <= 12'd1949;
            6'd32: Q <= 12'd873;
            6'd33: Q <= 12'd1630;
            6'd34: Q <= 12'd1936;
            6'd35: Q <= 12'd2624;
            6'd36: Q <= 12'd2798;
            6'd37: Q <= 12'd2063;
            6'd38: Q <= 12'd1568;
            6'd39: Q <= 12'd2529;
            6'd40: Q <= 12'd1664;
            6'd41: Q <= 12'd3309;
            6'd42: Q <= 12'd2039;
            6'd43: Q <= 12'd315;
            6'd44: Q <= 12'd2008;
            6'd45: Q <= 12'd424;
            6'd46: Q <= 12'd716;
            6'd47: Q <= 12'd987;
            6'd48: Q <= 12'd2075;
            6'd49: Q <= 12'd3104;
            6'd50: Q <= 12'd468;
            6'd51: Q <= 12'd1047;
            6'd52: Q <= 12'd2616;
            6'd53: Q <= 12'd1441;
            6'd54: Q <= 12'd1397;
            6'd55: Q <= 12'd2888;
            6'd56: Q <= 12'd3181;
            6'd57: Q <= 12'd738;
            6'd58: Q <= 12'd995;
            6'd59: Q <= 12'd28;
            6'd60: Q <= 12'd1806;
            6'd61: Q <= 12'd2331;
            6'd62: Q <= 12'd2209;
        endcase  
    end
    
endmodule
    
module tf1_ROM (
    input                       clk,
    input      [4:0]            A,
    output reg [23:0]           Q
);
    
    always@(posedge clk) begin
        case(A)
            5'd0: Q <= 24'b101111101100000110111011;
            5'd1: Q <= 24'b010000110011010001000101;
            5'd2: Q <= 24'b001000100010011110000111;
            5'd3: Q <= 24'b001000000001010110110111;
            5'd4: Q <= 24'b100000111011010000110101;
            5'd5: Q <= 24'b110000111100100011100010;
            5'd6: Q <= 24'b001001011110100110100100;
            5'd7: Q <= 24'b100010000011100101011000;
            5'd8: Q <= 24'b010011010001010100010001;
            5'd9: Q <= 24'b011110011001001001100111;
            5'd10: Q <= 24'b011100100000010001101101;
            5'd11: Q <= 24'b011111111011000100010110;
            5'd12: Q <= 24'b010001111101100111101001;
            5'd13: Q <= 24'b011001001010001010000110;
            5'd14: Q <= 24'b101101111011010111000101;
            5'd15: Q <= 24'b100110110111100011101100;
            5'd16: Q <= 24'b110001100100010111110101;
            5'd17: Q <= 24'b010000110110101110000111;
            5'd18: Q <= 24'b010100110011001111000000;
            5'd19: Q <= 24'b011011110101000000011000;
            5'd20: Q <= 24'b101111100101011001111000;
            5'd21: Q <= 24'b101110101101010101011101;
            5'd22: Q <= 24'b011111101010001101001110;
            5'd23: Q <= 24'b001000100110100010001001;
            5'd24: Q <= 24'b000010000110011111000001;
            5'd25: Q <= 24'b101100010001010100010010;
            5'd26: Q <= 24'b010010000010010010101011;
            5'd27: Q <= 24'b010010101010000110111110;
            5'd28: Q <= 24'b100110111010001100101101;
            5'd29: Q <= 24'b100111111111000100001110;
            5'd30: Q <= 24'b000111011100001011100101;
            5'd31: Q <= 24'b101111000000001110100110;
        endcase  
    end

endmodule

