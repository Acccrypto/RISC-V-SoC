// Actel Corporation Proprietary and Confidential
// Copyright 2008 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN 
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED 
// IN ADVANCE IN WRITING.  
// Revision Information:
// SVN Revision Information:
// SVN $Revision: 6419 $
// SVN $Date: 2009-02-04 04:34:22 -0800 (Wed, 04 Feb 2009) $
`timescale 1ns/100ps
module
GPIO_GPIO_0_BFM_MAIN // BFM_MAIN changed to BFM_MAIN_GPIO so that it should not take internal BFM.
(
SYSCLK
,
SYSRSTN
,
PCLK
,
HCLK
,
HRESETN
,
HADDR
,
HBURST
,
HMASTLOCK
,
HPROT
,
HSIZE
,
HTRANS
,
HWRITE
,
HWDATA
,
HRDATA
,
HREADY
,
HRESP
,
HSEL
,
INTERRUPT
,
GP_OUT
,
GP_IN
,
EXT_WR
,
EXT_RD
,
EXT_ADDR
,
EXT_DATA
,
EXT_WAIT
,
CON_ADDR
,
CON_DATA
,
CON_RD
,
CON_WR
,
CON_BUSY
,
INSTR_OUT
,
INSTR_IN
,
FINISHED
,
FAILED
)
;
parameter
OPMODE
=
0
;
parameter
VECTFILE
=
"test.vec"
;
parameter
MAX_INSTRUCTIONS
=
16384
;
parameter
MAX_STACK
=
1024
;
parameter
MAX_MEMTEST
=
65536
;
parameter
TPD
=
1
;
parameter
DEBUGLEVEL
=
-
1
;
parameter
CON_SPULSE
=
0
;
parameter
ARGVALUE0
=
0
;
parameter
ARGVALUE1
=
0
;
parameter
ARGVALUE2
=
0
;
parameter
ARGVALUE3
=
0
;
parameter
ARGVALUE4
=
0
;
parameter
ARGVALUE5
=
0
;
parameter
ARGVALUE6
=
0
;
parameter
ARGVALUE7
=
0
;
parameter
ARGVALUE8
=
0
;
parameter
ARGVALUE9
=
0
;
parameter
ARGVALUE10
=
0
;
parameter
ARGVALUE11
=
0
;
parameter
ARGVALUE12
=
0
;
parameter
ARGVALUE13
=
0
;
parameter
ARGVALUE14
=
0
;
parameter
ARGVALUE15
=
0
;
parameter
ARGVALUE16
=
0
;
parameter
ARGVALUE17
=
0
;
parameter
ARGVALUE18
=
0
;
parameter
ARGVALUE19
=
0
;
parameter
ARGVALUE20
=
0
;
parameter
ARGVALUE21
=
0
;
parameter
ARGVALUE22
=
0
;
parameter
ARGVALUE23
=
0
;
parameter
ARGVALUE24
=
0
;
parameter
ARGVALUE25
=
0
;
parameter
ARGVALUE26
=
0
;
parameter
ARGVALUE27
=
0
;
parameter
ARGVALUE28
=
0
;
parameter
ARGVALUE29
=
0
;
parameter
ARGVALUE30
=
0
;
parameter
ARGVALUE31
=
0
;
parameter
ARGVALUE32
=
0
;
parameter
ARGVALUE33
=
0
;
parameter
ARGVALUE34
=
0
;
parameter
ARGVALUE35
=
0
;
parameter
ARGVALUE36
=
0
;
parameter
ARGVALUE37
=
0
;
parameter
ARGVALUE38
=
0
;
parameter
ARGVALUE39
=
0
;
parameter
ARGVALUE40
=
0
;
parameter
ARGVALUE41
=
0
;
parameter
ARGVALUE42
=
0
;
parameter
ARGVALUE43
=
0
;
parameter
ARGVALUE44
=
0
;
parameter
ARGVALUE45
=
0
;
parameter
ARGVALUE46
=
0
;
parameter
ARGVALUE47
=
0
;
parameter
ARGVALUE48
=
0
;
parameter
ARGVALUE49
=
0
;
parameter
ARGVALUE50
=
0
;
parameter
ARGVALUE51
=
0
;
parameter
ARGVALUE52
=
0
;
parameter
ARGVALUE53
=
0
;
parameter
ARGVALUE54
=
0
;
parameter
ARGVALUE55
=
0
;
parameter
ARGVALUE56
=
0
;
parameter
ARGVALUE57
=
0
;
parameter
ARGVALUE58
=
0
;
parameter
ARGVALUE59
=
0
;
parameter
ARGVALUE60
=
0
;
parameter
ARGVALUE61
=
0
;
parameter
ARGVALUE62
=
0
;
parameter
ARGVALUE63
=
0
;
parameter
ARGVALUE64
=
0
;
parameter
ARGVALUE65
=
0
;
parameter
ARGVALUE66
=
0
;
parameter
ARGVALUE67
=
0
;
parameter
ARGVALUE68
=
0
;
parameter
ARGVALUE69
=
0
;
parameter
ARGVALUE70
=
0
;
parameter
ARGVALUE71
=
0
;
parameter
ARGVALUE72
=
0
;
parameter
ARGVALUE73
=
0
;
parameter
ARGVALUE74
=
0
;
parameter
ARGVALUE75
=
0
;
parameter
ARGVALUE76
=
0
;
parameter
ARGVALUE77
=
0
;
parameter
ARGVALUE78
=
0
;
parameter
ARGVALUE79
=
0
;
parameter
ARGVALUE80
=
0
;
parameter
ARGVALUE81
=
0
;
parameter
ARGVALUE82
=
0
;
parameter
ARGVALUE83
=
0
;
parameter
ARGVALUE84
=
0
;
parameter
ARGVALUE85
=
0
;
parameter
ARGVALUE86
=
0
;
parameter
ARGVALUE87
=
0
;
parameter
ARGVALUE88
=
0
;
parameter
ARGVALUE89
=
0
;
parameter
ARGVALUE90
=
0
;
parameter
ARGVALUE91
=
0
;
parameter
ARGVALUE92
=
0
;
parameter
ARGVALUE93
=
0
;
parameter
ARGVALUE94
=
0
;
parameter
ARGVALUE95
=
0
;
parameter
ARGVALUE96
=
0
;
parameter
ARGVALUE97
=
0
;
parameter
ARGVALUE98
=
0
;
parameter
ARGVALUE99
=
0
;
localparam
[
1
:
(
3
)
*
8
]
BFMA1O
=
"2.1"
;
localparam
[
1
:
(
7
)
*
8
]
BFMA1I
=
"22Dec08"
;
input
SYSCLK
;
input
SYSRSTN
;
output
PCLK
;
wire
PCLK
;
output
HCLK
;
wire
HCLK
;
output
HRESETN
;
wire
#
TPD
HRESETN
;
output
[
31
:
0
]
HADDR
;
wire
[
31
:
0
]
#
TPD
HADDR
;
output
[
2
:
0
]
HBURST
;
wire
[
2
:
0
]
#
TPD
HBURST
;
output
HMASTLOCK
;
wire
#
TPD
HMASTLOCK
;
output
[
3
:
0
]
HPROT
;
wire
[
3
:
0
]
#
TPD
HPROT
;
output
[
2
:
0
]
HSIZE
;
wire
[
2
:
0
]
#
TPD
HSIZE
;
output
[
1
:
0
]
HTRANS
;
wire
[
1
:
0
]
#
TPD
HTRANS
;
output
HWRITE
;
wire
#
TPD
HWRITE
;
output
[
31
:
0
]
HWDATA
;
wire
[
31
:
0
]
#
TPD
HWDATA
;
input
[
31
:
0
]
HRDATA
;
input
HREADY
;
input
HRESP
;
output
[
15
:
0
]
HSEL
;
wire
[
15
:
0
]
#
TPD
HSEL
;
input
[
255
:
0
]
INTERRUPT
;
output
[
31
:
0
]
GP_OUT
;
wire
[
31
:
0
]
#
TPD
GP_OUT
;
input
[
31
:
0
]
GP_IN
;
output
EXT_WR
;
wire
#
TPD
EXT_WR
;
output
EXT_RD
;
wire
#
TPD
EXT_RD
;
output
[
31
:
0
]
EXT_ADDR
;
wire
[
31
:
0
]
#
TPD
EXT_ADDR
;
inout
[
31
:
0
]
EXT_DATA
;
wire
[
31
:
0
]
#
TPD
EXT_DATA
;
input
EXT_WAIT
;
input
[
15
:
0
]
CON_ADDR
;
inout
[
31
:
0
]
CON_DATA
;
wire
[
31
:
0
]
#
TPD
CON_DATA
;
wire
[
31
:
0
]
BFMA1l
;
input
CON_RD
;
input
CON_WR
;
output
CON_BUSY
;
reg
CON_BUSY
;
output
[
31
:
0
]
INSTR_OUT
;
reg
[
31
:
0
]
INSTR_OUT
;
input
[
31
:
0
]
INSTR_IN
;
output
FINISHED
;
wire
#
TPD
FINISHED
;
output
FAILED
;
wire
#
TPD
FAILED
;
localparam
BFMA1OI
=
0
;
wire
BFMA1II
;
integer
BFMA1lI
[
0
:
255
]
;
integer
BFMA1Ol
[
0
:
MAX_INSTRUCTIONS
-
1
]
;
reg
BFMA1Il
;
reg
[
2
:
0
]
BFMA1ll
;
reg
BFMA1O0
;
reg
[
3
:
0
]
BFMA1I0
;
reg
[
1
:
0
]
BFMA1l0
;
reg
BFMA1O1
;
wire
[
31
:
0
]
BFMA1I1
;
reg
[
31
:
0
]
BFMA1l1
;
reg
[
31
:
0
]
BFMA1OOI
;
reg
[
2
:
0
]
BFMA1IOI
;
reg
[
2
:
0
]
BFMA1lOI
;
reg
[
15
:
0
]
BFMA1OII
;
reg
BFMA1III
;
reg
BFMA1lII
;
reg
BFMA1OlI
;
reg
BFMA1IlI
;
reg
BFMA1llI
;
reg
BFMA1O0I
;
reg
BFMA1I0I
;
reg
BFMA1l0I
;
reg
[
31
:
0
]
BFMA1O1I
;
reg
[
31
:
0
]
BFMA1I1I
;
reg
[
31
:
0
]
BFMA1l1I
;
reg
[
31
:
0
]
BFMA1OOl
;
reg
[
31
:
0
]
BFMA1IOl
;
reg
[
31
:
0
]
BFMA1lOl
;
reg
[
31
:
0
]
BFMA1OIl
;
reg
[
31
:
0
]
BFMA1IIl
;
integer
BFMA1lIl
;
reg
BFMA1Oll
;
reg
BFMA1Ill
;
reg
[
31
:
0
]
BFMA1lll
;
reg
[
31
:
0
]
BFMA1O0l
;
integer
BFMA1I0l
;
reg
BFMA1l0l
;
reg
BFMA1O1l
;
reg
BFMA1I1l
;
reg
BFMA1l1l
;
reg
BFMA1OO0
;
wire
[
31
:
0
]
BFMA1IO0
;
reg
[
31
:
0
]
BFMA1lO0
;
reg
[
31
:
0
]
BFMA1OI0
;
reg
[
31
:
0
]
BFMA1II0
;
wire
[
31
:
0
]
BFMA1lI0
;
reg
[
31
:
0
]
BFMA1Ol0
;
reg
BFMA1Il0
;
reg
BFMA1ll0
;
integer
BFMA1O00
;
integer
BFMA1I00
;
reg
BFMA1l00
=
1
'b
0
;
reg
[
31
:
0
]
BFMA1O10
;
reg
[
1
:
(
80
)
*
8
]
BFMA1I10
;
reg
BFMA1l10
;
reg
BFMA1OO1
;
reg
BFMA1IO1
;
reg
BFMA1lO1
;
reg
BFMA1OI1
;
reg
BFMA1II1
;
parameter
[
31
:
0
]
BFMA1lI1
=
{
32
{
1
'b
0
}
}
;
parameter
[
255
:
0
]
BFMA1Ol1
=
{
256
{
1
'b
0
}
}
;
parameter
BFMA1Il1
=
TPD
*
1
;
assign
BFMA1II
=
SYSCLK
;
integer
BFMA1ll1
[
0
:
MAX_STACK
-
1
]
;
integer
BFMA1O01
;
integer
BFMA1I01
;
integer
BFMA1l01
;
integer
DEBUG
;
integer
BFMA1O11
;
// Actel Corporation Proprietary and Confidential
// Copyright 2008 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN 
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED 
// IN ADVANCE IN WRITING.  
// Revision Information:
// SVN Revision Information:
// SVN $Revision: 6419 $
// SVN $Date: 2009-02-04 04:34:22 -0800 (Wed, 04 Feb 2009) $
localparam
BFMA1I11
=
22
;
localparam
BFMA1l11
=
0
;
localparam
BFMA1OOOI
=
4
;
localparam
BFMA1IOOI
=
8
;
localparam
BFMA1lOOI
=
12
;
localparam
BFMA1OIOI
=
16
;
localparam
BFMA1IIOI
=
20
;
localparam
BFMA1lIOI
=
24
;
localparam
BFMA1OlOI
=
28
;
localparam
BFMA1IlOI
=
32
;
localparam
BFMA1llOI
=
36
;
localparam
BFMA1O0OI
=
40
;
localparam
BFMA1I0OI
=
44
;
localparam
BFMA1l0OI
=
48
;
localparam
BFMA1O1OI
=
52
;
localparam
BFMA1I1OI
=
56
;
localparam
BFMA1l1OI
=
60
;
localparam
BFMA1OOII
=
64
;
localparam
BFMA1IOII
=
68
;
localparam
BFMA1lOII
=
72
;
localparam
BFMA1OIII
=
76
;
localparam
BFMA1IIII
=
80
;
localparam
BFMA1lIII
=
100
;
localparam
BFMA1OlII
=
101
;
localparam
BFMA1IlII
=
102
;
localparam
BFMA1llII
=
103
;
localparam
BFMA1O0II
=
104
;
localparam
BFMA1I0II
=
105
;
localparam
BFMA1l0II
=
106
;
localparam
BFMA1O1II
=
107
;
localparam
BFMA1I1II
=
108
;
localparam
BFMA1l1II
=
109
;
localparam
BFMA1OOlI
=
110
;
localparam
BFMA1IOlI
=
111
;
localparam
BFMA1lOlI
=
112
;
localparam
BFMA1OIlI
=
113
;
localparam
BFMA1IIlI
=
114
;
localparam
BFMA1lIlI
=
115
;
localparam
BFMA1OllI
=
128
;
localparam
BFMA1IllI
=
129
;
localparam
BFMA1lllI
=
130
;
localparam
BFMA1O0lI
=
131
;
localparam
BFMA1I0lI
=
132
;
localparam
BFMA1l0lI
=
133
;
localparam
BFMA1O1lI
=
134
;
localparam
BFMA1I1lI
=
135
;
localparam
BFMA1l1lI
=
136
;
localparam
BFMA1OO0I
=
137
;
localparam
BFMA1IO0I
=
138
;
localparam
BFMA1lO0I
=
139
;
localparam
BFMA1OI0I
=
140
;
localparam
BFMA1II0I
=
141
;
localparam
BFMA1lI0I
=
142
;
localparam
BFMA1Ol0I
=
150
;
localparam
BFMA1Il0I
=
151
;
localparam
BFMA1ll0I
=
152
;
localparam
BFMA1O00I
=
153
;
localparam
BFMA1I00I
=
154
;
localparam
BFMA1l00I
=
160
;
localparam
BFMA1O10I
=
161
;
localparam
BFMA1I10I
=
162
;
localparam
BFMA1l10I
=
163
;
localparam
BFMA1OO1I
=
164
;
localparam
BFMA1IO1I
=
165
;
localparam
BFMA1lO1I
=
166
;
localparam
BFMA1OI1I
=
167
;
localparam
BFMA1II1I
=
168
;
localparam
BFMA1lI1I
=
169
;
localparam
BFMA1Ol1I
=
170
;
localparam
BFMA1Il1I
=
171
;
localparam
BFMA1ll1I
=
172
;
localparam
BFMA1O01I
=
200
;
localparam
BFMA1I01I
=
201
;
localparam
BFMA1l01I
=
202
;
localparam
BFMA1O11I
=
203
;
localparam
BFMA1I11I
=
204
;
localparam
BFMA1l11I
=
205
;
localparam
BFMA1OOOl
=
206
;
localparam
BFMA1IOOl
=
207
;
localparam
BFMA1lOOl
=
208
;
localparam
BFMA1OIOl
=
209
;
localparam
BFMA1IIOl
=
210
;
localparam
BFMA1lIOl
=
211
;
localparam
BFMA1OlOl
=
212
;
localparam
BFMA1IlOl
=
213
;
localparam
BFMA1llOl
=
214
;
localparam
BFMA1O0Ol
=
215
;
localparam
BFMA1I0Ol
=
216
;
localparam
BFMA1l0Ol
=
217
;
localparam
BFMA1O1Ol
=
218
;
localparam
BFMA1I1Ol
=
219
;
localparam
BFMA1l1Ol
=
220
;
localparam
BFMA1OOIl
=
221
;
localparam
BFMA1IOIl
=
222
;
localparam
BFMA1lOIl
=
250
;
localparam
BFMA1OIIl
=
251
;
localparam
BFMA1IIIl
=
252
;
localparam
BFMA1lIIl
=
253
;
localparam
BFMA1OlIl
=
254
;
localparam
BFMA1IlIl
=
255
;
localparam
BFMA1llIl
=
1001
;
localparam
BFMA1O0Il
=
1002
;
localparam
BFMA1I0Il
=
1003
;
localparam
BFMA1l0Il
=
1004
;
localparam
BFMA1O1Il
=
1005
;
localparam
BFMA1I1Il
=
1006
;
localparam
BFMA1l1Il
=
1007
;
localparam
BFMA1OOll
=
1008
;
localparam
BFMA1IOll
=
1009
;
localparam
BFMA1lOll
=
1010
;
localparam
BFMA1OIll
=
1011
;
localparam
BFMA1IIll
=
1012
;
localparam
BFMA1lIll
=
1013
;
localparam
BFMA1Olll
=
1014
;
localparam
BFMA1Illl
=
1015
;
localparam
BFMA1llll
=
1016
;
localparam
BFMA1O0ll
=
1017
;
localparam
BFMA1I0ll
=
1018
;
localparam
BFMA1l0ll
=
1019
;
localparam
BFMA1O1ll
=
1020
;
localparam
BFMA1I1ll
=
1021
;
localparam
BFMA1l1ll
=
1022
;
localparam
BFMA1OO0l
=
1023
;
localparam
BFMA1IO0l
=
0
;
localparam
BFMA1lO0l
=
1
;
localparam
BFMA1OI0l
=
2
;
localparam
BFMA1II0l
=
3
;
localparam
BFMA1lI0l
=
4
;
localparam
BFMA1Ol0l
=
5
;
localparam
BFMA1Il0l
=
6
;
localparam
BFMA1ll0l
=
7
;
localparam
BFMA1O00l
=
8
;
localparam
BFMA1I00l
=
0
;
localparam
BFMA1l00l
=
1
;
localparam
BFMA1O10l
=
2
;
localparam
BFMA1I10l
=
3
;
localparam
BFMA1l10l
=
4
;
localparam
BFMA1OO1l
=
32
'h
00000000
;
localparam
BFMA1IO1l
=
32
'h
00002000
;
localparam
BFMA1lO1l
=
32
'h
00004000
;
localparam
BFMA1OI1l
=
32
'h
00006000
;
localparam
BFMA1II1l
=
32
'h
00008000
;
localparam
[
1
:
0
]
BFMA1lI1l
=
0
;
localparam
[
1
:
0
]
BFMA1Ol1l
=
1
;
localparam
[
1
:
0
]
BFMA1Il1l
=
2
;
localparam
[
1
:
0
]
BFMA1ll1l
=
3
;
function
integer
BFMA1O01l
;
input
[
31
:
0
]
BFMA1I01l
;
integer
BFMA1ll1l
;
begin
BFMA1ll1l
=
BFMA1I01l
;
BFMA1O01l
=
BFMA1ll1l
;
end
endfunction
function
integer
to_int_unsigned
;
input
[
31
:
0
]
BFMA1I01l
;
integer
BFMA1I01l
;
integer
BFMA1ll1l
;
begin
BFMA1ll1l
=
BFMA1I01l
;
to_int_unsigned
=
BFMA1ll1l
;
end
endfunction
function
integer
to_int_signed
;
input
[
31
:
0
]
BFMA1I01l
;
integer
BFMA1ll1l
;
begin
BFMA1ll1l
=
BFMA1I01l
;
to_int_signed
=
BFMA1ll1l
;
end
endfunction
function
[
31
:
0
]
to_slv32
;
input
BFMA1ll1l
;
integer
BFMA1ll1l
;
reg
[
31
:
0
]
BFMA1I01l
;
begin
BFMA1I01l
=
BFMA1ll1l
;
to_slv32
=
BFMA1I01l
;
end
endfunction
function
[
31
:
0
]
BFMA1l01l
;
input
[
2
:
0
]
BFMA1O11l
;
input
[
1
:
0
]
BFMA1I11l
;
input
[
31
:
0
]
BFMA1l11l
;
input
BFMA1OOO0
;
integer
BFMA1OOO0
;
reg
[
31
:
0
]
BFMA1IOO0
;
reg
BFMA1lOO0
;
begin
BFMA1IOO0
=
{
32
{
1
'b
0
}
}
;
case
(
BFMA1OOO0
)
0
:
begin
case
(
BFMA1O11l
)
3
'b
000
:
begin
case
(
BFMA1I11l
)
2
'b
00
:
begin
BFMA1IOO0
[
7
:
0
]
=
BFMA1l11l
[
7
:
0
]
;
end
2
'b
01
:
begin
BFMA1IOO0
[
15
:
8
]
=
BFMA1l11l
[
7
:
0
]
;
end
2
'b
10
:
begin
BFMA1IOO0
[
23
:
16
]
=
BFMA1l11l
[
7
:
0
]
;
end
2
'b
11
:
begin
BFMA1IOO0
[
31
:
24
]
=
BFMA1l11l
[
7
:
0
]
;
end
default
:
begin
end
endcase
end
3
'b
001
:
begin
case
(
BFMA1I11l
)
2
'b
00
:
begin
BFMA1IOO0
[
15
:
0
]
=
BFMA1l11l
[
15
:
0
]
;
end
2
'b
01
:
begin
BFMA1IOO0
[
15
:
0
]
=
BFMA1l11l
[
15
:
0
]
;
$display
(
"BFM: Missaligned AHB Cycle(Half A10=01) ? (WARNING)"
)
;
end
2
'b
10
:
begin
BFMA1IOO0
[
31
:
16
]
=
BFMA1l11l
[
15
:
0
]
;
end
2
'b
11
:
begin
BFMA1IOO0
[
31
:
16
]
=
BFMA1l11l
[
15
:
0
]
;
$display
(
"BFM: Missaligned AHB Cycle(Half A10=11) ? (WARNING)"
)
;
end
default
:
begin
end
endcase
end
3
'b
010
:
begin
BFMA1IOO0
=
BFMA1l11l
;
case
(
BFMA1I11l
)
2
'b
00
:
begin
end
2
'b
01
:
begin
$display
(
"BFM: Missaligned AHB Cycle(Word A10=01) ? (WARNING)"
)
;
end
2
'b
10
:
begin
$display
(
"BFM: Missaligned AHB Cycle(Word A10=10) ? (WARNING)"
)
;
end
2
'b
11
:
begin
$display
(
"BFM: Missaligned AHB Cycle(Word A10=11) ? (WARNING)"
)
;
end
default
:
begin
end
endcase
end
default
:
begin
$display
(
"Unexpected AHB Size setting (ERROR)"
)
;
end
endcase
end
1
:
begin
case
(
BFMA1O11l
)
3
'b
000
:
begin
case
(
BFMA1I11l
)
2
'b
00
:
begin
BFMA1IOO0
[
7
:
0
]
=
BFMA1l11l
[
7
:
0
]
;
end
2
'b
01
:
begin
BFMA1IOO0
[
15
:
8
]
=
BFMA1l11l
[
7
:
0
]
;
end
2
'b
10
:
begin
BFMA1IOO0
[
7
:
0
]
=
BFMA1l11l
[
7
:
0
]
;
end
2
'b
11
:
begin
BFMA1IOO0
[
15
:
8
]
=
BFMA1l11l
[
7
:
0
]
;
end
default
:
begin
end
endcase
end
3
'b
001
:
begin
BFMA1IOO0
[
15
:
0
]
=
BFMA1l11l
[
15
:
0
]
;
case
(
BFMA1I11l
)
2
'b
00
:
begin
end
2
'b
01
:
begin
$display
(
"BFM: Missaligned AHB Cycle(Half A10=01) ? (WARNING)"
)
;
end
2
'b
10
:
begin
$display
(
"BFM: Missaligned AHB Cycle(Half A10=10) ? (WARNING)"
)
;
end
2
'b
11
:
begin
$display
(
"BFM: Missaligned AHB Cycle(Half A10=11) ? (WARNING)"
)
;
end
default
:
begin
end
endcase
end
default
:
begin
$display
(
"Unexpected AHB Size setting (ERROR)"
)
;
end
endcase
end
2
:
begin
case
(
BFMA1O11l
)
3
'b
000
:
begin
BFMA1IOO0
[
7
:
0
]
=
BFMA1l11l
[
7
:
0
]
;
end
default
:
begin
$display
(
"Unexpected AHB Size setting (ERROR)"
)
;
end
endcase
end
8
:
begin
BFMA1IOO0
=
BFMA1l11l
;
end
default
:
begin
$display
(
"Illegal Alignment mode (ERROR)"
)
;
end
endcase
BFMA1l01l
=
BFMA1IOO0
;
end
endfunction
function
[
31
:
0
]
BFMA1OIO0
;
input
[
2
:
0
]
BFMA1O11l
;
input
[
1
:
0
]
BFMA1I11l
;
input
[
31
:
0
]
BFMA1l11l
;
input
BFMA1OOO0
;
integer
BFMA1OOO0
;
reg
[
31
:
0
]
BFMA1IOO0
;
begin
BFMA1IOO0
=
BFMA1l01l
(
BFMA1O11l
,
BFMA1I11l
,
BFMA1l11l
,
BFMA1OOO0
)
;
BFMA1OIO0
=
BFMA1IOO0
;
end
endfunction
function
[
31
:
0
]
BFMA1IIO0
;
input
[
2
:
0
]
BFMA1O11l
;
input
[
1
:
0
]
BFMA1I11l
;
input
[
31
:
0
]
BFMA1l11l
;
input
BFMA1OOO0
;
integer
BFMA1OOO0
;
reg
[
31
:
0
]
BFMA1IOO0
;
reg
BFMA1lOO0
;
begin
if
(
BFMA1OOO0
==
8
)
begin
BFMA1IOO0
=
BFMA1l11l
;
end
else
begin
BFMA1IOO0
=
0
;
BFMA1lOO0
=
BFMA1I11l
[
1
]
;
case
(
BFMA1O11l
)
3
'b
000
:
begin
case
(
BFMA1I11l
)
2
'b
00
:
BFMA1IOO0
[
7
:
0
]
=
BFMA1l11l
[
7
:
0
]
;
2
'b
01
:
BFMA1IOO0
[
7
:
0
]
=
BFMA1l11l
[
15
:
8
]
;
2
'b
10
:
BFMA1IOO0
[
7
:
0
]
=
BFMA1l11l
[
23
:
16
]
;
2
'b
11
:
BFMA1IOO0
[
7
:
0
]
=
BFMA1l11l
[
31
:
24
]
;
default
:
begin
end
endcase
end
3
'b
001
:
begin
case
(
BFMA1lOO0
)
1
'b
0
:
BFMA1IOO0
[
15
:
0
]
=
BFMA1l11l
[
15
:
0
]
;
1
'b
1
:
BFMA1IOO0
[
15
:
0
]
=
BFMA1l11l
[
31
:
16
]
;
default
:
begin
end
endcase
end
3
'b
010
:
begin
BFMA1IOO0
=
BFMA1l11l
;
end
default
:
$display
(
"Unexpected AHB Size setting (ERROR)"
)
;
endcase
end
BFMA1IIO0
=
BFMA1IOO0
;
end
endfunction
function
integer
BFMA1lIO0
;
input
BFMA1ll1l
;
integer
BFMA1ll1l
;
integer
BFMA1OlO0
;
begin
BFMA1OlO0
=
BFMA1ll1l
;
BFMA1lIO0
=
BFMA1OlO0
;
end
endfunction
function
integer
BFMA1IlO0
;
input
BFMA1O11l
;
integer
BFMA1O11l
;
integer
BFMA1OlO0
;
begin
case
(
BFMA1O11l
)
0
:
begin
BFMA1OlO0
=
'h
62
;
end
1
:
begin
BFMA1OlO0
=
'h
68
;
end
2
:
begin
BFMA1OlO0
=
'h
77
;
end
3
:
begin
BFMA1OlO0
=
'h
78
;
end
default
:
begin
BFMA1OlO0
=
'h
3f
;
end
endcase
BFMA1IlO0
=
BFMA1OlO0
;
end
endfunction
function
integer
BFMA1llO0
;
input
BFMA1O11l
;
integer
BFMA1O11l
;
input
BFMA1O0O0
;
integer
BFMA1O0O0
;
integer
BFMA1OlO0
;
begin
case
(
BFMA1O11l
)
0
:
begin
BFMA1OlO0
=
1
;
end
1
:
begin
BFMA1OlO0
=
2
;
end
2
:
begin
BFMA1OlO0
=
4
;
end
3
:
begin
BFMA1OlO0
=
BFMA1O0O0
;
end
default
:
begin
BFMA1OlO0
=
0
;
end
endcase
BFMA1llO0
=
BFMA1OlO0
;
end
endfunction
function
integer
BFMA1I0O0
;
input
BFMA1O11l
;
integer
BFMA1O11l
;
input
BFMA1l0O0
;
integer
BFMA1l0O0
;
reg
[
2
:
0
]
BFMA1OlO0
;
begin
case
(
BFMA1O11l
)
0
:
begin
BFMA1OlO0
=
3
'b
000
;
end
1
:
begin
BFMA1OlO0
=
3
'b
001
;
end
2
:
begin
BFMA1OlO0
=
3
'b
010
;
end
3
:
begin
BFMA1OlO0
=
BFMA1l0O0
;
end
default
:
begin
BFMA1OlO0
=
3
'b
XXX
;
end
endcase
BFMA1I0O0
=
BFMA1OlO0
;
end
endfunction
function
integer
BFMA1O1O0
;
input
BFMA1I1O0
;
integer
BFMA1I1O0
;
input
BFMA1ll1l
;
integer
BFMA1ll1l
;
input
BFMA1l1O0
;
integer
BFMA1l1O0
;
input
BFMA1OOI0
;
integer
BFMA1OOI0
;
integer
BFMA1IOI0
;
reg
[
31
:
0
]
BFMA1lOI0
;
reg
[
31
:
0
]
BFMA1OII0
;
reg
[
31
:
0
]
BFMA1III0
;
integer
BFMA1lII0
;
reg
[
63
:
0
]
BFMA1OlI0
;
localparam
[
31
:
0
]
BFMA1IlI0
=
0
;
localparam
[
31
:
0
]
BFMA1llI0
=
1
;
begin
BFMA1lOI0
=
BFMA1ll1l
;
BFMA1OII0
=
BFMA1l1O0
;
BFMA1lII0
=
BFMA1l1O0
;
BFMA1III0
=
{
32
{
1
'b
0
}
}
;
case
(
BFMA1I1O0
)
BFMA1llIl
:
begin
BFMA1III0
=
0
;
end
BFMA1O0Il
:
begin
BFMA1III0
=
BFMA1lOI0
+
BFMA1OII0
;
end
BFMA1I0Il
:
begin
BFMA1III0
=
BFMA1lOI0
-
BFMA1OII0
;
end
BFMA1l0Il
:
begin
BFMA1OlI0
=
BFMA1lOI0
*
BFMA1OII0
;
BFMA1III0
=
BFMA1OlI0
[
31
:
0
]
;
end
BFMA1O1Il
:
begin
BFMA1III0
=
BFMA1lOI0
/
BFMA1OII0
;
end
BFMA1OOll
:
begin
BFMA1III0
=
BFMA1lOI0
&
BFMA1OII0
;
end
BFMA1IOll
:
begin
BFMA1III0
=
BFMA1lOI0
|
BFMA1OII0
;
end
BFMA1lOll
:
begin
BFMA1III0
=
BFMA1lOI0
^
BFMA1OII0
;
end
BFMA1OIll
:
begin
BFMA1III0
=
BFMA1lOI0
^
BFMA1OII0
;
end
BFMA1lIll
:
begin
if
(
BFMA1lII0
==
0
)
begin
BFMA1III0
=
BFMA1lOI0
;
end
else
begin
BFMA1III0
=
BFMA1lOI0
>>
BFMA1lII0
;
end
end
BFMA1IIll
:
begin
if
(
BFMA1lII0
==
0
)
begin
BFMA1III0
=
BFMA1lOI0
;
end
else
begin
BFMA1III0
=
BFMA1lOI0
<<
BFMA1lII0
;
end
end
BFMA1l1Il
:
begin
BFMA1OlI0
=
{
BFMA1IlI0
,
BFMA1llI0
}
;
if
(
BFMA1lII0
>
0
)
begin
begin
:
BFMA1O0I0
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
1
;
BFMA1I0I0
<=
BFMA1lII0
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
BFMA1OlI0
=
BFMA1OlI0
[
31
:
0
]
*
BFMA1lOI0
;
end
end
end
BFMA1III0
=
BFMA1OlI0
[
31
:
0
]
;
end
BFMA1Olll
:
begin
if
(
BFMA1lOI0
==
BFMA1OII0
)
begin
BFMA1III0
=
BFMA1llI0
;
end
end
BFMA1Illl
:
begin
if
(
BFMA1lOI0
!=
BFMA1OII0
)
begin
BFMA1III0
=
BFMA1llI0
;
end
end
BFMA1llll
:
begin
if
(
BFMA1lOI0
>
BFMA1OII0
)
begin
BFMA1III0
=
BFMA1llI0
;
end
end
BFMA1O0ll
:
begin
if
(
BFMA1lOI0
<
BFMA1OII0
)
begin
BFMA1III0
=
BFMA1llI0
;
end
end
BFMA1I0ll
:
begin
if
(
BFMA1lOI0
>=
BFMA1OII0
)
begin
BFMA1III0
=
BFMA1llI0
;
end
end
BFMA1l0ll
:
begin
if
(
BFMA1lOI0
<=
BFMA1OII0
)
begin
BFMA1III0
=
BFMA1llI0
;
end
end
BFMA1I1Il
:
begin
BFMA1III0
=
BFMA1lOI0
%
BFMA1OII0
;
end
BFMA1O1ll
:
begin
if
(
BFMA1l1O0
<=
31
)
begin
BFMA1III0
=
BFMA1lOI0
;
BFMA1III0
[
BFMA1l1O0
]
=
1
'b
1
;
end
else
begin
$display
(
"Bit operation on bit >31 (FAILURE)"
)
;
$stop
;
end
end
BFMA1I1ll
:
begin
if
(
BFMA1l1O0
<=
31
)
begin
BFMA1III0
=
BFMA1lOI0
;
BFMA1III0
[
BFMA1l1O0
]
=
1
'b
0
;
end
else
begin
$display
(
"Bit operation on bit >31 (FAILURE)"
)
;
$stop
;
end
end
BFMA1l1ll
:
begin
if
(
BFMA1l1O0
<=
31
)
begin
BFMA1III0
=
BFMA1lOI0
;
BFMA1III0
[
BFMA1l1O0
]
=
~
BFMA1III0
[
BFMA1l1O0
]
;
end
else
begin
$display
(
"Bit operation on bit >31 (FAILURE)"
)
;
$stop
;
end
end
BFMA1OO0l
:
begin
if
(
BFMA1l1O0
<=
31
)
begin
BFMA1III0
=
0
;
BFMA1III0
[
0
]
=
BFMA1lOI0
[
BFMA1l1O0
]
;
end
else
begin
$display
(
"Bit operation on bit >31 (FAILURE)"
)
;
$stop
;
end
end
default
:
begin
$display
(
"Illegal Maths Operator (FAILURE)"
)
;
$stop
;
end
endcase
BFMA1IOI0
=
BFMA1III0
;
if
(
BFMA1OOI0
>=
4
)
begin
$display
(
"Calculated %d = %d (%d) %d"
,
BFMA1IOI0
,
BFMA1ll1l
,
BFMA1I1O0
,
BFMA1l1O0
)
;
end
BFMA1O1O0
=
BFMA1IOI0
;
end
endfunction
function
[
31
:
0
]
BFMA1l0I0
;
input
[
31
:
0
]
BFMA1ll1l
;
reg
[
31
:
0
]
BFMA1O1I0
;
begin
BFMA1O1I0
=
BFMA1ll1l
;
BFMA1O1I0
=
0
;
begin
:
BFMA1I1I0
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
31
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
if
(
(
BFMA1ll1l
[
BFMA1I0I0
]
)
==
1
'b
1
)
begin
BFMA1O1I0
[
BFMA1I0I0
]
=
1
'b
1
;
end
end
end
BFMA1l0I0
=
BFMA1O1I0
;
end
endfunction
function
integer
BFMA1l1I0
;
input
BFMA1OOl0
;
integer
BFMA1OOl0
;
input
BFMA1ll1l
;
integer
BFMA1ll1l
;
integer
BFMA1IOl0
;
integer
BFMA1lOl0
;
begin
BFMA1lOl0
=
BFMA1OOl0
/
BFMA1ll1l
;
BFMA1IOl0
=
BFMA1OOl0
-
BFMA1lOl0
*
BFMA1ll1l
;
BFMA1l1I0
=
BFMA1IOl0
;
end
endfunction
function
integer
BFMA1OIl0
;
input
BFMA1OOl0
;
integer
BFMA1OOl0
;
input
BFMA1ll1l
;
integer
BFMA1ll1l
;
integer
BFMA1IOl0
;
integer
BFMA1lOl0
;
begin
BFMA1lOl0
=
BFMA1OOl0
/
BFMA1ll1l
;
BFMA1IOl0
=
BFMA1OOl0
-
BFMA1lOl0
*
BFMA1ll1l
;
BFMA1OIl0
=
BFMA1lOl0
;
end
endfunction
function
integer
to_boolean
;
input
BFMA1ll1l
;
integer
BFMA1ll1l
;
integer
BFMA1IIl0
;
begin
BFMA1IIl0
=
0
;
if
(
BFMA1ll1l
!=
0
)
BFMA1IIl0
=
1
;
to_boolean
=
BFMA1IIl0
;
end
endfunction
function
integer
BFMA1lIl0
;
input
BFMA1Oll0
;
integer
BFMA1Oll0
;
reg
[
31
:
0
]
BFMA1Ill0
;
reg
[
31
:
0
]
BFMA1lll0
;
reg
BFMA1O0l0
;
begin
BFMA1Ill0
=
BFMA1Oll0
;
BFMA1O0l0
=
1
'b
1
;
BFMA1lll0
[
0
]
=
BFMA1O0l0
^
BFMA1Ill0
[
31
]
;
BFMA1lll0
[
1
]
=
BFMA1O0l0
^
BFMA1Ill0
[
31
]
^
BFMA1Ill0
[
0
]
;
BFMA1lll0
[
2
]
=
BFMA1O0l0
^
BFMA1Ill0
[
31
]
^
BFMA1Ill0
[
1
]
;
BFMA1lll0
[
3
]
=
BFMA1Ill0
[
2
]
;
BFMA1lll0
[
4
]
=
BFMA1O0l0
^
BFMA1Ill0
[
31
]
^
BFMA1Ill0
[
3
]
;
BFMA1lll0
[
5
]
=
BFMA1O0l0
^
BFMA1Ill0
[
31
]
^
BFMA1Ill0
[
4
]
;
BFMA1lll0
[
6
]
=
BFMA1Ill0
[
5
]
;
BFMA1lll0
[
7
]
=
BFMA1O0l0
^
BFMA1Ill0
[
31
]
^
BFMA1Ill0
[
6
]
;
BFMA1lll0
[
8
]
=
BFMA1O0l0
^
BFMA1Ill0
[
31
]
^
BFMA1Ill0
[
7
]
;
BFMA1lll0
[
9
]
=
BFMA1Ill0
[
8
]
;
BFMA1lll0
[
10
]
=
BFMA1O0l0
^
BFMA1Ill0
[
31
]
^
BFMA1Ill0
[
9
]
;
BFMA1lll0
[
11
]
=
BFMA1O0l0
^
BFMA1Ill0
[
31
]
^
BFMA1Ill0
[
10
]
;
BFMA1lll0
[
12
]
=
BFMA1O0l0
^
BFMA1Ill0
[
31
]
^
BFMA1Ill0
[
11
]
;
BFMA1lll0
[
13
]
=
BFMA1Ill0
[
12
]
;
BFMA1lll0
[
14
]
=
BFMA1Ill0
[
13
]
;
BFMA1lll0
[
15
]
=
BFMA1Ill0
[
14
]
;
BFMA1lll0
[
16
]
=
BFMA1O0l0
^
BFMA1Ill0
[
31
]
^
BFMA1Ill0
[
15
]
;
BFMA1lll0
[
17
]
=
BFMA1Ill0
[
16
]
;
BFMA1lll0
[
18
]
=
BFMA1Ill0
[
17
]
;
BFMA1lll0
[
19
]
=
BFMA1Ill0
[
18
]
;
BFMA1lll0
[
20
]
=
BFMA1Ill0
[
19
]
;
BFMA1lll0
[
21
]
=
BFMA1Ill0
[
20
]
;
BFMA1lll0
[
22
]
=
BFMA1O0l0
^
BFMA1Ill0
[
31
]
^
BFMA1Ill0
[
21
]
;
BFMA1lll0
[
23
]
=
BFMA1O0l0
^
BFMA1Ill0
[
31
]
^
BFMA1Ill0
[
22
]
;
BFMA1lll0
[
24
]
=
BFMA1Ill0
[
23
]
;
BFMA1lll0
[
25
]
=
BFMA1Ill0
[
24
]
;
BFMA1lll0
[
26
]
=
BFMA1O0l0
^
BFMA1Ill0
[
31
]
^
BFMA1Ill0
[
25
]
;
BFMA1lll0
[
27
]
=
BFMA1Ill0
[
26
]
;
BFMA1lll0
[
28
]
=
BFMA1Ill0
[
27
]
;
BFMA1lll0
[
29
]
=
BFMA1Ill0
[
28
]
;
BFMA1lll0
[
30
]
=
BFMA1Ill0
[
29
]
;
BFMA1lll0
[
31
]
=
BFMA1Ill0
[
30
]
;
BFMA1lIl0
=
BFMA1lll0
;
end
endfunction
function
integer
BFMA1I0l0
;
input
BFMA1Oll0
;
integer
BFMA1Oll0
;
input
BFMA1O11l
;
integer
BFMA1O11l
;
integer
BFMA1l0l0
;
integer
BFMA1I0I0
;
reg
[
31
:
0
]
BFMA1Ill0
;
begin
BFMA1Ill0
=
BFMA1Oll0
;
for
(
BFMA1I0I0
=
31
;
BFMA1I0I0
>=
BFMA1O11l
;
BFMA1I0I0
=
BFMA1I0I0
-
1
)
BFMA1Ill0
[
BFMA1I0I0
]
=
0
;
BFMA1l0l0
=
BFMA1Ill0
;
BFMA1I0l0
=
BFMA1l0l0
;
end
endfunction
function
integer
BFMA1O1l0
;
input
BFMA1Oll0
;
integer
BFMA1Oll0
;
input
BFMA1O11l
;
integer
BFMA1O11l
;
integer
BFMA1l0l0
;
reg
[
31
:
0
]
BFMA1Ill0
;
integer
BFMA1I1l0
;
integer
BFMA1I0I0
;
begin
case
(
BFMA1O11l
)
1
:
begin
BFMA1I1l0
=
0
;
end
2
:
begin
BFMA1I1l0
=
1
;
end
4
:
begin
BFMA1I1l0
=
2
;
end
8
:
begin
BFMA1I1l0
=
3
;
end
16
:
begin
BFMA1I1l0
=
4
;
end
32
:
begin
BFMA1I1l0
=
5
;
end
64
:
begin
BFMA1I1l0
=
6
;
end
128
:
begin
BFMA1I1l0
=
7
;
end
256
:
begin
BFMA1I1l0
=
8
;
end
512
:
begin
BFMA1I1l0
=
9
;
end
1024
:
begin
BFMA1I1l0
=
10
;
end
2048
:
begin
BFMA1I1l0
=
11
;
end
4096
:
begin
BFMA1I1l0
=
12
;
end
8192
:
begin
BFMA1I1l0
=
13
;
end
16384
:
begin
BFMA1I1l0
=
14
;
end
32768
:
begin
BFMA1I1l0
=
15
;
end
65536
:
begin
BFMA1I1l0
=
16
;
end
131072
:
BFMA1I1l0
=
17
;
262144
:
BFMA1I1l0
=
18
;
524288
:
BFMA1I1l0
=
19
;
1048576
:
BFMA1I1l0
=
20
;
2097152
:
BFMA1I1l0
=
21
;
4194304
:
BFMA1I1l0
=
22
;
8388608
:
BFMA1I1l0
=
23
;
16777216
:
BFMA1I1l0
=
24
;
33554432
:
BFMA1I1l0
=
25
;
67108864
:
BFMA1I1l0
=
26
;
134217728
:
BFMA1I1l0
=
27
;
268435456
:
BFMA1I1l0
=
28
;
536870912
:
BFMA1I1l0
=
29
;
1073741824
:
BFMA1I1l0
=
30
;
default
:
begin
$display
(
"Random function error (FAILURE)"
)
;
$finish
;
end
endcase
BFMA1Ill0
=
to_slv32
(
BFMA1Oll0
)
;
if
(
BFMA1I1l0
<
31
)
begin
for
(
BFMA1I0I0
=
31
;
BFMA1I0I0
>=
BFMA1I1l0
;
BFMA1I0I0
=
BFMA1I0I0
-
1
)
BFMA1Ill0
[
BFMA1I0I0
]
=
0
;
end
BFMA1l0l0
=
to_int_signed
(
BFMA1Ill0
)
;
BFMA1O1l0
=
BFMA1l0l0
;
end
endfunction
function
bound1k
;
input
BFMA1l1l0
;
integer
BFMA1l1l0
;
input
BFMA1OO00
;
integer
BFMA1OO00
;
reg
[
31
:
0
]
BFMA1IO00
;
reg
BFMA1lO00
;
begin
BFMA1IO00
=
BFMA1OO00
;
BFMA1lO00
=
0
;
case
(
BFMA1l1l0
)
0
:
begin
if
(
BFMA1IO00
[
9
:
0
]
==
10
'b
0000000000
)
begin
BFMA1lO00
=
1
;
end
end
1
:
begin
BFMA1lO00
=
1
;
end
2
:
begin
end
default
:
begin
$display
(
"Illegal Burst Boundary Set (FAILURE)"
)
;
$finish
;
end
endcase
bound1k
=
BFMA1lO00
;
end
endfunction
function
integer
BFMA1OI00
;
input
BFMA1II00
;
integer
BFMA1II00
;
integer
BFMA1lI00
;
integer
BFMA1Ol00
;
integer
BFMA1Il00
;
begin
BFMA1Ol00
=
BFMA1II00
/
65536
;
BFMA1lI00
=
BFMA1II00
%
65536
;
BFMA1Il00
=
2
+
BFMA1lI00
+
1
+
(
(
BFMA1Ol00
-
1
)
/
4
)
;
BFMA1OI00
=
BFMA1Il00
;
end
endfunction
function
[
1
:
(
256
)
*
8
]
BFMA1ll00
;
input
BFMA1O000
;
integer
BFMA1O000
;
reg
[
1
:
(
256
)
*
8
]
BFMA1I000
;
reg
[
1
:
(
256
)
*
8
]
BFMA1l000
;
integer
BFMA1I0I0
;
integer
BFMA1O100
;
integer
BFMA1I100
;
reg
[
31
:
0
]
BFMA1l100
;
integer
BFMA1lI00
;
integer
BFMA1Ol00
;
integer
BFMA1II00
;
integer
BFMA1OO10
;
begin
BFMA1Ol00
=
BFMA1Ol
[
BFMA1O000
+
1
]
/
65536
;
BFMA1lI00
=
BFMA1Ol
[
BFMA1O000
+
1
]
%
65536
;
BFMA1II00
=
2
+
BFMA1lI00
+
1
+
(
(
BFMA1Ol00
-
1
)
/
4
)
;
for
(
BFMA1O100
=
1
;
BFMA1O100
<=
256
*
8
;
BFMA1O100
=
BFMA1O100
+
1
)
BFMA1I000
[
BFMA1O100
]
=
0
;
BFMA1I0I0
=
BFMA1O000
+
2
+
BFMA1lI00
;
BFMA1I100
=
3
;
begin
:
BFMA1IO10
integer
BFMA1O100
;
for
(
BFMA1O100
=
1
;
BFMA1O100
<=
BFMA1Ol00
;
BFMA1O100
=
BFMA1O100
+
1
)
begin
BFMA1l100
=
BFMA1Ol
[
BFMA1I0I0
]
;
for
(
BFMA1OO10
=
1
;
BFMA1OO10
<=
8
;
BFMA1OO10
=
BFMA1OO10
+
1
)
BFMA1I000
[
(
BFMA1O100
-
1
)
*
8
+
BFMA1OO10
]
=
BFMA1l100
[
BFMA1I100
*
8
+
8
-
BFMA1OO10
]
;
if
(
BFMA1I100
==
0
)
begin
BFMA1I0I0
=
BFMA1I0I0
+
1
;
BFMA1I100
=
4
;
end
BFMA1I100
=
BFMA1I100
-
1
;
end
end
case
(
BFMA1lI00
)
0
:
begin
$sformat
(
BFMA1l000
,
BFMA1I000
)
;
end
1
:
begin
$sformat
(
BFMA1l000
,
BFMA1I000
,
BFMA1lI
[
2
]
)
;
end
2
:
begin
$sformat
(
BFMA1l000
,
BFMA1I000
,
BFMA1lI
[
2
]
,
BFMA1lI
[
3
]
)
;
end
3
:
begin
$sformat
(
BFMA1l000
,
BFMA1I000
,
BFMA1lI
[
2
]
,
BFMA1lI
[
3
]
,
BFMA1lI
[
4
]
)
;
end
4
:
begin
$sformat
(
BFMA1l000
,
BFMA1I000
,
BFMA1lI
[
2
]
,
BFMA1lI
[
3
]
,
BFMA1lI
[
4
]
,
BFMA1lI
[
5
]
)
;
end
5
:
begin
$sformat
(
BFMA1l000
,
BFMA1I000
,
BFMA1lI
[
2
]
,
BFMA1lI
[
3
]
,
BFMA1lI
[
4
]
,
BFMA1lI
[
5
]
,
BFMA1lI
[
6
]
)
;
end
6
:
begin
$sformat
(
BFMA1l000
,
BFMA1I000
,
BFMA1lI
[
2
]
,
BFMA1lI
[
3
]
,
BFMA1lI
[
4
]
,
BFMA1lI
[
5
]
,
BFMA1lI
[
6
]
,
BFMA1lI
[
7
]
)
;
end
7
:
begin
$sformat
(
BFMA1l000
,
BFMA1I000
,
BFMA1lI
[
2
]
,
BFMA1lI
[
3
]
,
BFMA1lI
[
4
]
,
BFMA1lI
[
5
]
,
BFMA1lI
[
6
]
,
BFMA1lI
[
7
]
,
BFMA1lI
[
8
]
)
;
end
default
:
begin
$display
(
"String Error (FAILURE)"
)
;
end
endcase
BFMA1ll00
=
BFMA1l000
;
end
endfunction
integer
BFMA1lO10
;
integer
BFMA1OI10
;
integer
BFMA1II10
;
integer
BFMA1lI10
;
parameter
[
2
:
0
]
BFMA1Ol10
=
0
;
parameter
[
2
:
0
]
BFMA1Il10
=
1
;
parameter
[
2
:
0
]
BFMA1ll10
=
2
;
parameter
[
2
:
0
]
BFMA1O010
=
3
;
parameter
[
2
:
0
]
BFMA1I010
=
4
;
parameter
[
2
:
0
]
BFMA1l010
=
5
;
integer
BFMA1O110
;
integer
BFMA1I110
;
integer
BFMA1l110
;
integer
BFMA1OOO1
;
integer
BFMA1IOO1
;
reg
[
2
:
0
]
BFMA1lOO1
;
integer
BFMA1OIO1
[
0
:
MAX_MEMTEST
-
1
]
;
integer
BFMA1IIO1
;
integer
BFMA1lIO1
;
integer
BFMA1OlO1
;
integer
BFMA1IlO1
;
reg
BFMA1llO1
;
integer
BFMA1O0O1
;
integer
BFMA1I0O1
;
integer
BFMA1l0O1
;
integer
BFMA1O1O1
;
integer
BFMA1I1O1
;
integer
BFMA1l1O1
;
reg
BFMA1OOI1
;
reg
BFMA1IOI1
;
reg
BFMA1lOI1
;
reg
BFMA1OII1
;
integer
BFMA1III1
;
function
automatic
integer
BFMA1lII1
;
input
BFMA1OlI1
;
input
BFMA1IlI1
;
integer
BFMA1IlI1
;
integer
BFMA1llI1
;
integer
BFMA1O0I1
;
integer
BFMA1I0I1
;
integer
BFMA1l0I1
;
integer
BFMA1O1I1
;
integer
BFMA1I1I1
;
reg
[
31
:
0
]
BFMA1I01l
;
integer
BFMA1l1I1
;
begin
if
(
BFMA1OlI1
)
begin
BFMA1I01l
=
BFMA1IlI1
;
BFMA1O0I1
=
BFMA1I01l
[
30
:
16
]
;
BFMA1I0I1
=
BFMA1I01l
[
14
:
13
]
;
BFMA1l0I1
=
BFMA1I01l
[
12
:
0
]
;
BFMA1O1I1
=
BFMA1I01l
[
12
:
8
]
;
BFMA1I1I1
=
BFMA1I01l
[
7
:
0
]
;
BFMA1l1I1
=
0
;
if
(
(
BFMA1I01l
[
15
]
)
==
1
'b
1
)
begin
BFMA1l1I1
=
BFMA1lII1
(
1
,
BFMA1O0I1
)
;
end
case
(
BFMA1I0I1
)
3
:
begin
case
(
BFMA1O1I1
)
BFMA1I00l
:
begin
case
(
BFMA1I1I1
)
BFMA1lO0l
:
begin
BFMA1llI1
=
BFMA1O01
;
end
BFMA1OI0l
:
begin
BFMA1llI1
=
(
$time
/
1
)
;
end
BFMA1II0l
:
begin
BFMA1llI1
=
DEBUG
;
end
BFMA1lI0l
:
begin
BFMA1llI1
=
BFMA1l01
;
end
BFMA1Ol0l
:
begin
BFMA1llI1
=
BFMA1II10
;
end
BFMA1Il0l
:
begin
BFMA1llI1
=
BFMA1l1O1
-
1
;
end
BFMA1ll0l
:
begin
BFMA1llI1
=
BFMA1O1O1
;
end
BFMA1O00l
:
begin
BFMA1llI1
=
BFMA1I1O1
;
end
default
:
begin
$display
(
"Illegal Parameter P0 (FAILURE)"
)
;
end
endcase
end
BFMA1l00l
:
begin
case
(
BFMA1I1I1
)
0
:
BFMA1llI1
=
ARGVALUE0
;
1
:
BFMA1llI1
=
ARGVALUE1
;
2
:
BFMA1llI1
=
ARGVALUE2
;
3
:
BFMA1llI1
=
ARGVALUE3
;
4
:
BFMA1llI1
=
ARGVALUE4
;
5
:
BFMA1llI1
=
ARGVALUE5
;
6
:
BFMA1llI1
=
ARGVALUE6
;
7
:
BFMA1llI1
=
ARGVALUE7
;
8
:
BFMA1llI1
=
ARGVALUE8
;
9
:
BFMA1llI1
=
ARGVALUE9
;
10
:
BFMA1llI1
=
ARGVALUE10
;
11
:
BFMA1llI1
=
ARGVALUE11
;
12
:
BFMA1llI1
=
ARGVALUE12
;
13
:
BFMA1llI1
=
ARGVALUE13
;
14
:
BFMA1llI1
=
ARGVALUE14
;
15
:
BFMA1llI1
=
ARGVALUE15
;
16
:
BFMA1llI1
=
ARGVALUE16
;
17
:
BFMA1llI1
=
ARGVALUE17
;
18
:
BFMA1llI1
=
ARGVALUE18
;
19
:
BFMA1llI1
=
ARGVALUE19
;
20
:
BFMA1llI1
=
ARGVALUE20
;
21
:
BFMA1llI1
=
ARGVALUE21
;
22
:
BFMA1llI1
=
ARGVALUE22
;
23
:
BFMA1llI1
=
ARGVALUE23
;
24
:
BFMA1llI1
=
ARGVALUE24
;
25
:
BFMA1llI1
=
ARGVALUE25
;
26
:
BFMA1llI1
=
ARGVALUE26
;
27
:
BFMA1llI1
=
ARGVALUE27
;
28
:
BFMA1llI1
=
ARGVALUE28
;
29
:
BFMA1llI1
=
ARGVALUE29
;
30
:
BFMA1llI1
=
ARGVALUE30
;
31
:
BFMA1llI1
=
ARGVALUE31
;
32
:
BFMA1llI1
=
ARGVALUE32
;
33
:
BFMA1llI1
=
ARGVALUE33
;
34
:
BFMA1llI1
=
ARGVALUE34
;
35
:
BFMA1llI1
=
ARGVALUE35
;
36
:
BFMA1llI1
=
ARGVALUE36
;
37
:
BFMA1llI1
=
ARGVALUE37
;
38
:
BFMA1llI1
=
ARGVALUE38
;
39
:
BFMA1llI1
=
ARGVALUE39
;
40
:
BFMA1llI1
=
ARGVALUE40
;
41
:
BFMA1llI1
=
ARGVALUE41
;
42
:
BFMA1llI1
=
ARGVALUE42
;
43
:
BFMA1llI1
=
ARGVALUE43
;
44
:
BFMA1llI1
=
ARGVALUE44
;
45
:
BFMA1llI1
=
ARGVALUE45
;
46
:
BFMA1llI1
=
ARGVALUE46
;
47
:
BFMA1llI1
=
ARGVALUE47
;
48
:
BFMA1llI1
=
ARGVALUE48
;
49
:
BFMA1llI1
=
ARGVALUE49
;
50
:
BFMA1llI1
=
ARGVALUE50
;
51
:
BFMA1llI1
=
ARGVALUE51
;
52
:
BFMA1llI1
=
ARGVALUE52
;
53
:
BFMA1llI1
=
ARGVALUE53
;
54
:
BFMA1llI1
=
ARGVALUE54
;
55
:
BFMA1llI1
=
ARGVALUE55
;
56
:
BFMA1llI1
=
ARGVALUE56
;
57
:
BFMA1llI1
=
ARGVALUE57
;
58
:
BFMA1llI1
=
ARGVALUE58
;
59
:
BFMA1llI1
=
ARGVALUE59
;
60
:
BFMA1llI1
=
ARGVALUE60
;
61
:
BFMA1llI1
=
ARGVALUE61
;
62
:
BFMA1llI1
=
ARGVALUE62
;
63
:
BFMA1llI1
=
ARGVALUE63
;
64
:
BFMA1llI1
=
ARGVALUE64
;
65
:
BFMA1llI1
=
ARGVALUE65
;
66
:
BFMA1llI1
=
ARGVALUE66
;
67
:
BFMA1llI1
=
ARGVALUE67
;
68
:
BFMA1llI1
=
ARGVALUE68
;
69
:
BFMA1llI1
=
ARGVALUE69
;
70
:
BFMA1llI1
=
ARGVALUE70
;
71
:
BFMA1llI1
=
ARGVALUE71
;
72
:
BFMA1llI1
=
ARGVALUE72
;
73
:
BFMA1llI1
=
ARGVALUE73
;
74
:
BFMA1llI1
=
ARGVALUE74
;
75
:
BFMA1llI1
=
ARGVALUE75
;
76
:
BFMA1llI1
=
ARGVALUE76
;
77
:
BFMA1llI1
=
ARGVALUE77
;
78
:
BFMA1llI1
=
ARGVALUE78
;
79
:
BFMA1llI1
=
ARGVALUE79
;
80
:
BFMA1llI1
=
ARGVALUE80
;
81
:
BFMA1llI1
=
ARGVALUE81
;
82
:
BFMA1llI1
=
ARGVALUE82
;
83
:
BFMA1llI1
=
ARGVALUE83
;
84
:
BFMA1llI1
=
ARGVALUE84
;
85
:
BFMA1llI1
=
ARGVALUE85
;
86
:
BFMA1llI1
=
ARGVALUE86
;
87
:
BFMA1llI1
=
ARGVALUE87
;
88
:
BFMA1llI1
=
ARGVALUE88
;
89
:
BFMA1llI1
=
ARGVALUE89
;
90
:
BFMA1llI1
=
ARGVALUE90
;
91
:
BFMA1llI1
=
ARGVALUE91
;
92
:
BFMA1llI1
=
ARGVALUE92
;
93
:
BFMA1llI1
=
ARGVALUE93
;
94
:
BFMA1llI1
=
ARGVALUE94
;
95
:
BFMA1llI1
=
ARGVALUE95
;
96
:
BFMA1llI1
=
ARGVALUE96
;
97
:
BFMA1llI1
=
ARGVALUE97
;
98
:
BFMA1llI1
=
ARGVALUE98
;
99
:
BFMA1llI1
=
ARGVALUE99
;
default
:
begin
$display
(
"Illegal Parameter P1 (FAILURE)"
)
;
end
endcase
end
BFMA1O10l
:
begin
BFMA1lO10
=
BFMA1lIl0
(
BFMA1lO10
)
;
BFMA1llI1
=
BFMA1I0l0
(
BFMA1lO10
,
BFMA1I1I1
)
;
end
BFMA1I10l
:
begin
BFMA1OI10
=
BFMA1lO10
;
BFMA1lO10
=
BFMA1lIl0
(
BFMA1lO10
)
;
BFMA1llI1
=
BFMA1I0l0
(
BFMA1lO10
,
BFMA1I1I1
)
;
end
BFMA1l10l
:
begin
BFMA1lO10
=
BFMA1OI10
;
BFMA1lO10
=
BFMA1lIl0
(
BFMA1lO10
)
;
BFMA1llI1
=
BFMA1I0l0
(
BFMA1lO10
,
BFMA1I1I1
)
;
end
default
:
begin
$display
(
"Illegal Parameter P2 (FAILURE)"
)
;
end
endcase
end
2
:
begin
BFMA1llI1
=
BFMA1ll1
[
BFMA1I01
-
BFMA1l0I1
+
BFMA1l1I1
]
;
end
1
:
begin
BFMA1llI1
=
BFMA1ll1
[
BFMA1l0I1
+
BFMA1l1I1
]
;
end
0
:
begin
BFMA1llI1
=
BFMA1l0I1
;
end
default
:
begin
$display
(
"Illegal Parameter P3 (FAILURE)"
)
;
end
endcase
end
else
begin
BFMA1llI1
=
BFMA1IlI1
;
end
BFMA1lII1
=
BFMA1llI1
;
end
endfunction
function
integer
BFMA1OOl1
;
input
BFMA1IlI1
;
integer
BFMA1IlI1
;
input
BFMA1I01
;
integer
BFMA1I01
;
integer
BFMA1IOl1
;
integer
BFMA1O0I1
;
integer
BFMA1I0I1
;
integer
BFMA1l0I1
;
integer
BFMA1O1I1
;
integer
BFMA1I1I1
;
reg
[
31
:
0
]
BFMA1I01l
;
integer
BFMA1l1I1
;
begin
BFMA1I01l
=
BFMA1IlI1
;
BFMA1O0I1
=
BFMA1I01l
[
30
:
16
]
;
BFMA1I0I1
=
BFMA1I01l
[
14
:
13
]
;
BFMA1l0I1
=
BFMA1I01l
[
12
:
0
]
;
BFMA1O1I1
=
BFMA1I01l
[
12
:
8
]
;
BFMA1I1I1
=
BFMA1I01l
[
7
:
0
]
;
BFMA1l1I1
=
0
;
if
(
(
BFMA1I01l
[
15
]
)
==
1
'b
1
)
begin
BFMA1l1I1
=
BFMA1lII1
(
1
,
BFMA1O0I1
)
;
end
case
(
BFMA1I0I1
)
3
:
begin
$display
(
"$Variables not allowed (FAILURE)"
)
;
end
2
:
begin
BFMA1IOl1
=
BFMA1I01
-
BFMA1l0I1
+
BFMA1l1I1
;
end
1
:
begin
BFMA1IOl1
=
BFMA1l0I1
+
BFMA1l1I1
;
end
0
:
begin
$display
(
"Immediate data not allowed (FAILURE)"
)
;
end
default
:
begin
$display
(
"Illegal Parameter P3 (FAILURE)"
)
;
end
endcase
BFMA1OOl1
=
BFMA1IOl1
;
end
endfunction
always
@
(
posedge
BFMA1II
or
negedge
SYSRSTN
)
begin
:
BFMA1lOl1
parameter
[
0
:
0
]
BFMA1OIl1
=
0
;
parameter
[
0
:
0
]
BFMA1IIl1
=
1
;
integer
BFMA1lIl1
;
reg
BFMA1Oll1
;
integer
BFMA1Ill1
[
0
:
4
]
;
reg
[
31
:
0
]
BFMA1lll1
[
0
:
255
]
;
integer
BFMA1O0l1
;
integer
BFMA1O000
;
integer
BFMA1I0l1
;
integer
BFMA1l0l1
;
integer
BFMA1O1l1
;
reg
[
31
:
0
]
BFMA1I1l1
;
reg
[
1
:
0
]
BFMA1l1l1
;
integer
BFMA1OO01
;
integer
BFMA1IO01
;
integer
BFMA1lO01
;
integer
BFMA1OI01
;
integer
BFMA1II01
;
reg
[
2
:
0
]
BFMA1lI01
;
reg
[
31
:
0
]
BFMA1Ol01
;
reg
[
31
:
0
]
BFMA1Il01
;
reg
[
31
:
0
]
BFMA1ll01
;
reg
BFMA1O001
;
reg
BFMA1I001
;
reg
BFMA1l001
;
reg
BFMA1O101
;
reg
BFMA1I101
;
reg
BFMA1l101
;
reg
BFMA1OO11
;
reg
BFMA1IO11
;
reg
BFMA1lO11
;
reg
BFMA1OI11
;
reg
BFMA1II11
;
integer
BFMA1lI11
;
integer
BFMA1Ol11
;
integer
BFMA1Il11
;
integer
BFMA1Il00
;
integer
BFMA1I0I0
;
integer
BFMA1I100
;
integer
BFMA1IlI1
;
integer
BFMA1llI1
;
integer
BFMA1ll11
;
reg
[
1
:
(
256
)
*
8
]
BFMA1l000
;
reg
[
1
:
(
256
)
*
8
]
BFMA1O011
;
reg
[
1
:
(
256
)
*
8
]
BFMA1I011
;
integer
BFMA1l011
;
integer
BFMA1O111
;
integer
BFMA1I111
;
integer
BFMA1l111
;
integer
BFMA1OOOOI
[
0
:
8191
]
;
reg
[
1
:
(
8
)
*
8
]
BFMA1IOOOI
;
reg
BFMA1lOOOI
;
reg
BFMA1OIOOI
;
reg
BFMA1IIOOI
;
integer
BFMA1lIOOI
;
integer
BFMA1OlOOI
;
integer
BFMA1IlOOI
;
integer
BFMA1llOOI
;
integer
BFMA1O0OOI
;
integer
BFMA1I0OOI
;
integer
BFMA1lI00
;
integer
BFMA1l0OOI
;
integer
BFMA1O1OOI
;
integer
BFMA1I1OOI
;
integer
BFMA1l1OOI
;
integer
BFMA1OOIOI
;
integer
BFMA1IOIOI
;
integer
BFMA1lOIOI
;
integer
BFMA1OIIOI
;
reg
[
31
:
0
]
BFMA1IIIOI
;
reg
[
31
:
0
]
BFMA1lIIOI
;
reg
BFMA1OlIOI
;
reg
BFMA1IlIOI
;
reg
BFMA1llIOI
;
reg
BFMA1O0IOI
;
reg
[
0
:
0
]
BFMA1I0IOI
;
reg
[
1
:
(
10
)
*
8
]
BFMA1l0IOI
;
reg
BFMA1O1IOI
;
reg
[
3
:
0
]
BFMA1I1IOI
;
reg
[
2
:
0
]
BFMA1l1IOI
;
integer
BFMA1OOlOI
;
reg
BFMA1IOlOI
;
reg
[
1
:
(
256
)
*
8
]
BFMA1lOlOI
[
0
:
100
]
;
integer
BFMA1OIlOI
;
integer
BFMA1IIlOI
;
reg
[
1
:
0
]
BFMA1lIlOI
;
reg
[
5
:
0
]
BFMA1OllOI
;
reg
[
16
:
0
]
BFMA1IllOI
;
reg
BFMA1lllOI
;
integer
BFMA1O0lOI
;
reg
BFMA1I0lOI
;
reg
BFMA1l0lOI
;
reg
BFMA1O1lOI
;
reg
BFMA1I1lOI
;
reg
BFMA1l1lOI
;
integer
BFMA1OO0OI
;
reg
BFMA1IO0OI
;
reg
BFMA1lO0OI
;
reg
BFMA1OI0OI
;
reg
BFMA1II0OI
;
reg
BFMA1lI0OI
;
integer
BFMA1Ol0OI
;
integer
BFMA1Il0OI
;
integer
BFMA1ll0OI
;
integer
BFMA1O00OI
;
reg
BFMA1I00OI
;
reg
[
1
:
0
]
BFMA1l00OI
;
reg
[
3
:
0
]
BFMA1O10OI
;
reg
[
2
:
0
]
BFMA1I10OI
;
reg
BFMA1l10OI
;
reg
BFMA1OO1OI
;
reg
[
256
*
8
:
0
]
BFMA1IO1OI
;
integer
BFMA1OlO0
;
integer
BFMA1OO10
;
integer
BFMA1lO1OI
;
reg
BFMA1OI1OI
;
integer
BFMA1OOI1
;
integer
BFMA1II1OI
[
0
:
15
]
;
integer
BFMA1lI1OI
;
integer
BFMA1Ol1OI
[
0
:
255
]
;
reg
[
8
:
0
]
BFMA1Il1OI
;
reg
[
8
:
0
]
BFMA1ll1OI
;
integer
BFMA1O01OI
[
0
:
255
]
;
integer
BFMA1I01OI
;
if
(
SYSRSTN
==
1
'b
0
)
begin
BFMA1OOIOI
=
0
;
BFMA1IOIOI
=
0
;
BFMA1II10
=
0
;
BFMA1OIlOI
=
0
;
BFMA1IIlOI
=
65536
;
BFMA1I0IOI
=
BFMA1OIl1
;
BFMA1lI10
=
0
;
BFMA1O1O1
=
0
;
BFMA1I1O1
=
0
;
BFMA1l00
<=
1
'b
0
;
DEBUG
<=
DEBUGLEVEL
;
BFMA1l1
<=
{
32
{
1
'b
0
}
}
;
BFMA1ll
<=
{
3
{
1
'b
0
}
}
;
BFMA1O0
<=
1
'b
0
;
BFMA1I0
<=
{
4
{
1
'b
0
}
}
;
BFMA1IOI
<=
{
3
{
1
'b
0
}
}
;
BFMA1l0
<=
{
2
{
1
'b
0
}
}
;
BFMA1O1
<=
1
'b
0
;
BFMA1O10
<=
{
32
{
1
'b
0
}
}
;
INSTR_OUT
<=
{
32
{
1
'b
0
}
}
;
BFMA1lII
<=
1
'b
0
;
BFMA1OlI
<=
1
'b
0
;
BFMA1O1I
<=
{
32
{
1
'b
0
}
}
;
BFMA1I1I
<=
{
32
{
1
'b
0
}
}
;
BFMA1l1I
<=
{
32
{
1
'b
0
}
}
;
BFMA1l1l
<=
1
'b
0
;
BFMA1l0l
<=
1
'b
0
;
BFMA1O1l
<=
1
'b
0
;
BFMA1OI0
<=
{
32
{
1
'b
0
}
}
;
BFMA1lO0
<=
{
32
{
1
'b
0
}
}
;
BFMA1l10
<=
1
'b
0
;
BFMA1I10
[
1
:
8
]
<=
{
"UNKNOWN"
,
8
'b
0
}
;
BFMA1IlI
<=
1
'b
0
;
BFMA1OOl
<=
{
32
{
1
'b
0
}
}
;
BFMA1IOl
<=
{
32
{
1
'b
0
}
}
;
BFMA1I00
<=
0
;
BFMA1OOI
<=
{
32
{
1
'b
0
}
}
;
BFMA1OO1
<=
1
'b
0
;
BFMA1Il
<=
1
'b
0
;
CON_BUSY
<=
1
'b
0
;
BFMA1I00
<=
0
;
BFMA1llI
<=
1
'b
0
;
BFMA1O0I
<=
1
'b
0
;
BFMA1IO1
<=
0
;
BFMA1lO1
<=
0
;
BFMA1OI1
<=
0
;
BFMA1II1
<=
0
;
BFMA1Oll1
=
0
;
BFMA1O000
=
0
;
BFMA1OI11
=
0
;
BFMA1l1OOI
=
0
;
BFMA1O001
=
0
;
BFMA1OO11
=
0
;
BFMA1I101
=
0
;
BFMA1I001
=
0
;
BFMA1l001
=
0
;
BFMA1O101
=
0
;
BFMA1l101
=
0
;
BFMA1IO11
=
0
;
BFMA1I01
=
0
;
BFMA1I1OOI
=
0
;
BFMA1II01
=
512
;
BFMA1IOlOI
=
0
;
BFMA1II10
=
0
;
BFMA1O0IOI
=
0
;
BFMA1O1IOI
=
1
'b
0
;
BFMA1I1IOI
=
4
'b
0011
;
BFMA1l1IOI
=
3
'b
001
;
BFMA1lOOOI
=
0
;
BFMA1lIlOI
=
2
;
BFMA1OllOI
=
4
;
BFMA1IllOI
=
0
;
BFMA1lllOI
=
0
;
BFMA1I0lOI
=
0
;
BFMA1l1lOI
=
0
;
BFMA1O01
=
0
;
BFMA1l0lOI
=
0
;
BFMA1OO0OI
=
0
;
BFMA1lO0OI
=
0
;
BFMA1OI0OI
=
0
;
BFMA1II0OI
=
0
;
BFMA1lI0OI
=
0
;
BFMA1O11
=
BFMA1OI
;
BFMA1IO0OI
=
0
;
BFMA1O00OI
=
0
;
BFMA1lO10
=
1
;
BFMA1OI10
=
1
;
BFMA1O11
=
1
;
BFMA1lI1OI
=
0
;
BFMA1Il1OI
=
0
;
BFMA1ll1OI
=
0
;
BFMA1I01OI
=
0
;
BFMA1O0lOI
=
0
;
end
else
begin
BFMA1Il0
<=
CON_RD
;
BFMA1ll0
<=
CON_WR
;
BFMA1l0l
<=
1
'b
0
;
BFMA1O1l
<=
1
'b
0
;
BFMA1l1l
<=
1
'b
0
;
BFMA1OO0
<=
1
'b
0
;
BFMA1lO11
=
0
;
if
(
~
BFMA1Oll1
)
begin
$display
(
" "
)
;
$display
(
"###########################################################################"
)
;
$display
(
"AMBA BFM Model"
)
;
$display
(
"Version %s %s"
,
BFMA1O
,
BFMA1I
)
;
$display
(
" "
)
;
$display
(
"Opening BFM Script file %0s"
,
VECTFILE
)
;
if
(
~
BFMA1Oll1
&
OPMODE
!=
2
)
begin
$readmemh
(
VECTFILE
,
BFMA1Ol
)
;
BFMA1ll11
=
3000
;
BFMA1Oll1
=
1
;
BFMA1O0l1
=
BFMA1Ol
[
4
]
;
BFMA1Ol0OI
=
BFMA1Ol
[
0
]
%
65536
;
BFMA1ll0OI
=
BFMA1Ol
[
0
]
/
65536
;
$display
(
"Read %0d Vectors - Compiler Version %0d.%0d"
,
BFMA1O0l1
,
BFMA1ll0OI
,
BFMA1Ol0OI
)
;
if
(
BFMA1ll0OI
!=
BFMA1I11
)
begin
$display
(
"Incorrect vectors file format for this BFM %0s  (FAILURE) == "
,
VECTFILE
)
;
$stop
;
end
BFMA1O000
=
BFMA1Ol
[
1
]
;
BFMA1l0l1
=
BFMA1Ol
[
2
]
;
BFMA1I01
=
BFMA1Ol
[
3
]
;
BFMA1ll1
[
BFMA1I01
]
=
0
;
BFMA1I01
=
BFMA1I01
+
1
;
if
(
BFMA1O000
==
0
)
begin
$display
(
"BFM Compiler reported errors (FAILURE)"
)
;
$stop
;
end
$display
(
"BFM:Filenames referenced in Vectors"
)
;
BFMA1I1l1
=
BFMA1Ol
[
BFMA1l0l1
]
;
BFMA1OO01
=
BFMA1Ol
[
BFMA1l0l1
]
%
256
;
while
(
BFMA1OO01
==
BFMA1ll0I
)
begin
BFMA1OI01
=
BFMA1OI00
(
BFMA1Ol
[
BFMA1l0l1
+
1
]
)
;
BFMA1l000
=
BFMA1ll00
(
BFMA1l0l1
)
;
$display
(
"  %0s"
,
BFMA1l000
)
;
begin
:
BFMA1l01OI
integer
BFMA1I0I0
,
BFMA1OO10
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<
256
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
for
(
BFMA1OO10
=
1
;
BFMA1OO10
<=
8
;
BFMA1OO10
=
BFMA1OO10
+
1
)
BFMA1lOlOI
[
BFMA1OIlOI
]
[
BFMA1I0I0
*
8
+
BFMA1OO10
]
=
BFMA1l000
[
BFMA1I0I0
*
8
+
BFMA1OO10
]
;
end
BFMA1OIlOI
=
BFMA1OIlOI
+
1
;
BFMA1l0l1
=
BFMA1l0l1
+
BFMA1OI01
;
BFMA1I1l1
=
to_slv32
(
BFMA1Ol
[
BFMA1l0l1
]
)
;
BFMA1OO01
=
BFMA1Ol
[
BFMA1l0l1
]
%
256
;
end
BFMA1IIlOI
=
65536
;
if
(
BFMA1OIlOI
>
1
)
BFMA1IIlOI
=
32768
;
if
(
BFMA1OIlOI
>
2
)
BFMA1IIlOI
=
16384
;
if
(
BFMA1OIlOI
>
4
)
BFMA1IIlOI
=
8912
;
if
(
BFMA1OIlOI
>
8
)
BFMA1IIlOI
=
4096
;
if
(
BFMA1OIlOI
>
16
)
BFMA1IIlOI
=
2048
;
if
(
BFMA1OIlOI
>
32
)
BFMA1IIlOI
=
1024
;
BFMA1l0lOI
=
(
OPMODE
==
0
)
;
end
end
if
(
OPMODE
==
2
&
~
BFMA1Oll1
)
begin
BFMA1IIlOI
=
65536
;
BFMA1Oll1
=
1
;
BFMA1l0lOI
=
0
;
BFMA1I01
=
BFMA1Ol
[
3
]
+
1
;
BFMA1ll1
[
BFMA1I01
]
=
0
;
BFMA1I01
=
BFMA1I01
+
1
;
end
if
(
BFMA1lI10
<=
1
)
begin
BFMA1Il
<=
1
'b
1
;
end
else
begin
BFMA1lI10
=
BFMA1lI10
-
1
;
end
case
(
BFMA1I0IOI
)
BFMA1OIl1
:
begin
if
(
HRESP
==
1
'b
1
&
HREADY
==
1
'b
1
)
begin
$display
(
"BFM: HRESP Signaling Protocol Error T2 (ERROR)"
)
;
BFMA1II10
=
BFMA1II10
+
1
;
end
if
(
HRESP
==
1
'b
1
&
HREADY
==
1
'b
0
)
begin
BFMA1I0IOI
=
BFMA1IIl1
;
end
end
BFMA1IIl1
:
begin
if
(
HRESP
==
1
'b
0
|
HREADY
==
1
'b
0
)
begin
$display
(
"BFM: HRESP Signaling Protocol Error T3 (ERROR)"
)
;
BFMA1II10
=
BFMA1II10
+
1
;
end
if
(
HRESP
==
1
'b
1
&
HREADY
==
1
'b
1
)
begin
BFMA1I0IOI
=
BFMA1OIl1
;
end
case
(
BFMA1I1OOI
)
0
:
begin
$display
(
"BFM: Unexpected HRESP Signaling Occured (ERROR)"
)
;
BFMA1II10
=
BFMA1II10
+
1
;
end
1
:
begin
BFMA1O0IOI
=
1
;
end
default
:
begin
$display
(
"BFM: HRESP mode is not correctly set (ERROR)"
)
;
BFMA1II10
=
BFMA1II10
+
1
;
end
endcase
end
endcase
if
(
OPMODE
>
0
)
begin
if
(
(
CON_WR
==
1
'b
1
)
&&
(
BFMA1ll0
==
1
'b
0
||
CON_SPULSE
==
1
)
)
begin
BFMA1Il00
=
BFMA1O01l
(
CON_ADDR
)
;
case
(
BFMA1Il00
)
0
:
begin
BFMA1l0lOI
=
(
(
BFMA1lI0
[
0
]
)
==
1
'b
1
)
;
BFMA1O1lOI
=
(
(
BFMA1lI0
[
1
]
)
==
1
'b
1
)
;
BFMA1lOOOI
=
0
;
if
(
BFMA1l0lOI
&
~
BFMA1O1lOI
)
begin
BFMA1ll1
[
BFMA1I01
]
=
0
;
BFMA1I01
=
BFMA1I01
+
1
;
end
if
(
DEBUG
>=
2
&
BFMA1l0lOI
&
~
BFMA1O1lOI
)
begin
$display
(
"BFM: Starting script at %08x (%0d parameters)"
,
BFMA1O000
,
BFMA1lI1OI
)
;
end
if
(
DEBUG
>=
2
&
BFMA1l0lOI
&
BFMA1O1lOI
)
begin
$display
(
"BFM: Starting instruction at %08x"
,
BFMA1O000
)
;
end
if
(
BFMA1l0lOI
)
begin
if
(
BFMA1lI1OI
>
0
)
begin
begin
:
BFMA1O11OI
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
BFMA1lI1OI
-
1
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
BFMA1ll1
[
BFMA1I01
]
=
BFMA1II1OI
[
BFMA1I0I0
]
;
BFMA1I01
=
BFMA1I01
+
1
;
end
end
BFMA1lI1OI
=
0
;
end
BFMA1Il1OI
=
0
;
BFMA1ll1OI
=
0
;
end
end
1
:
begin
BFMA1O000
=
BFMA1lI0
;
end
2
:
begin
BFMA1II1OI
[
BFMA1lI1OI
]
=
BFMA1lI0
;
BFMA1lI1OI
=
BFMA1lI1OI
+
1
;
end
default
:
begin
BFMA1Ol
[
BFMA1Il00
]
=
to_int_signed
(
BFMA1lI0
)
;
end
endcase
end
if
(
(
CON_RD
==
1
'b
1
)
&&
(
BFMA1Il0
==
1
'b
0
||
CON_SPULSE
==
1
)
)
begin
BFMA1Il00
=
BFMA1O01l
(
CON_ADDR
)
;
case
(
BFMA1Il00
)
0
:
begin
BFMA1Ol0
<=
{
32
{
1
'b
0
}
}
;
BFMA1Ol0
[
2
]
<=
BFMA1l0lOI
;
BFMA1Ol0
[
3
]
<=
(
BFMA1II10
>
0
)
;
end
1
:
begin
BFMA1Ol0
<=
BFMA1O000
;
end
2
:
begin
BFMA1Ol0
<=
BFMA1O01
;
BFMA1lI1OI
=
0
;
end
3
:
begin
if
(
BFMA1Il1OI
>
BFMA1ll1OI
)
begin
BFMA1Ol0
<=
BFMA1Ol1OI
[
BFMA1ll1OI
]
;
BFMA1ll1OI
=
BFMA1ll1OI
+
1
;
end
else
begin
$display
(
"BFM: Overread Control return stack"
)
;
BFMA1Ol0
<=
{
32
{
1
'b
0
}
}
;
end
end
default
:
begin
BFMA1Ol0
<=
{
32
{
1
'b
0
}
}
;
end
endcase
end
end
BFMA1OOIOI
=
BFMA1OOIOI
+
1
;
BFMA1l1O1
=
BFMA1l1O1
+
1
;
BFMA1OI1OI
=
1
;
while
(
BFMA1OI1OI
)
begin
BFMA1OI1OI
=
0
;
if
(
~
BFMA1OI11
&
BFMA1l0lOI
)
begin
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
7
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
BFMA1lI
[
BFMA1I0I0
]
=
0
;
BFMA1I1l1
=
BFMA1Ol
[
BFMA1O000
]
;
BFMA1l1l1
=
BFMA1I1l1
[
1
:
0
]
;
BFMA1OO01
=
BFMA1I1l1
[
7
:
0
]
;
BFMA1lO01
=
BFMA1I1l1
[
15
:
8
]
;
BFMA1l01
=
BFMA1I1l1
[
31
:
16
]
;
BFMA1Il11
=
BFMA1II01
;
BFMA1IOIOI
=
BFMA1IOIOI
+
1
;
BFMA1OI01
=
1
;
BFMA1OOlOI
=
-
1
;
BFMA1OO0OI
=
0
;
if
(
DEBUG
>=
5
)
$display
(
"BFM: Instruction %0d Line Number %0d Command %0d"
,
BFMA1O000
,
BFMA1l01
,
BFMA1OO01
)
;
if
(
BFMA1lI0OI
)
begin
$fdisplay
(
BFMA1lIl1
,
"%05d BF %4d %4d %3d"
,
$time
,
BFMA1O000
,
BFMA1l01
,
BFMA1OO01
)
;
end
if
(
BFMA1OO01
>=
100
)
begin
BFMA1IO01
=
BFMA1OO01
;
end
else
begin
BFMA1IO01
=
4
*
(
BFMA1OO01
/
4
)
;
end
if
(
BFMA1OO01
!=
BFMA1OI1I
)
begin
BFMA1OOIOI
=
0
;
end
case
(
BFMA1IO01
)
BFMA1Ol0I
,
BFMA1Il0I
,
BFMA1ll0I
,
BFMA1OIIl
:
BFMA1Il00
=
8
;
BFMA1IlOI
,
BFMA1l0OI
:
BFMA1Il00
=
4
+
BFMA1Ol
[
BFMA1O000
+
1
]
;
BFMA1l0lI
:
BFMA1Il00
=
3
+
BFMA1Ol
[
BFMA1O000
+
2
]
;
BFMA1I0lI
:
BFMA1Il00
=
3
;
BFMA1II0I
:
BFMA1Il00
=
2
+
BFMA1Ol
[
BFMA1O000
+
1
]
;
BFMA1I11I
:
BFMA1Il00
=
3
+
BFMA1Ol
[
BFMA1O000
+
2
]
;
BFMA1OlIl
:
BFMA1Il00
=
2
+
BFMA1Ol
[
BFMA1O000
+
1
]
;
BFMA1lIlI
:
BFMA1Il00
=
3
+
BFMA1Ol
[
BFMA1O000
+
1
]
;
default
:
BFMA1Il00
=
8
;
endcase
if
(
BFMA1Il00
>
0
)
begin
begin
:
BFMA1I11OI
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
BFMA1Il00
-
1
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
if
(
BFMA1I0I0
>=
1
&
BFMA1I0I0
<=
8
)
begin
BFMA1lI
[
BFMA1I0I0
]
=
BFMA1lII1
(
(
(
BFMA1I1l1
[
7
+
BFMA1I0I0
]
)
==
1
'b
1
)
,
BFMA1Ol
[
BFMA1O000
+
BFMA1I0I0
]
)
;
end
else
begin
BFMA1lI
[
BFMA1I0I0
]
=
BFMA1Ol
[
BFMA1O000
+
BFMA1I0I0
]
;
end
BFMA1lll1
[
BFMA1I0I0
]
=
to_slv32
(
BFMA1lI
[
BFMA1I0I0
]
)
;
end
end
end
case
(
BFMA1IO01
)
BFMA1IlIl
:
begin
$display
(
"BFM Compiler reported an error (FAILURE)"
)
;
BFMA1II10
=
BFMA1II10
+
1
;
$stop
;
end
BFMA1ll1I
:
begin
BFMA1OI01
=
2
;
BFMA1OI1OI
=
1
;
BFMA1Ol1OI
[
BFMA1Il1OI
]
=
BFMA1lI
[
1
]
;
BFMA1Il1OI
=
BFMA1Il1OI
+
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:conifpush %0d"
,
BFMA1l01
,
BFMA1lI
[
1
]
)
;
end
BFMA1OOOl
:
begin
BFMA1OI01
=
2
;
BFMA1Il
<=
1
'b
0
;
BFMA1lI10
=
BFMA1lI
[
1
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:RESET %0d"
,
BFMA1l01
,
BFMA1lI10
)
;
end
BFMA1IOOl
:
begin
BFMA1OI01
=
2
;
BFMA1l00
<=
BFMA1lll1
[
1
]
[
0
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:STOPCLK %0d "
,
BFMA1l01
,
BFMA1lll1
[
1
]
[
0
]
)
;
end
BFMA1l00I
:
begin
BFMA1OI01
=
2
;
BFMA1l1OOI
=
BFMA1lI
[
1
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:mode %0d (No effect in this version)"
,
BFMA1l01
,
BFMA1l1OOI
)
;
end
BFMA1O10I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
4
;
BFMA1Il00
=
BFMA1lI
[
1
]
;
BFMA1IlI1
=
BFMA1lI
[
2
]
;
BFMA1llI1
=
BFMA1lI
[
3
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:setup %0d %0d %0d "
,
BFMA1l01
,
BFMA1Il00
,
BFMA1IlI1
,
BFMA1llI1
)
;
case
(
BFMA1Il00
)
1
:
begin
BFMA1OI01
=
4
;
BFMA1lIlOI
=
BFMA1IlI1
;
BFMA1OllOI
=
BFMA1llI1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:Setup- Memory Cycle Transfer Size %0s %0d"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1lIlOI
)
,
BFMA1OllOI
)
;
end
2
:
begin
BFMA1OI01
=
3
;
BFMA1lllOI
=
to_boolean
(
BFMA1IlI1
)
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:Setup- Automatic Flush %0d"
,
BFMA1l01
,
BFMA1lllOI
)
;
end
3
:
begin
BFMA1OI01
=
3
;
BFMA1IllOI
=
BFMA1IlI1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:Setup- XRATE %0d"
,
BFMA1l01
,
BFMA1IllOI
)
;
end
4
:
begin
BFMA1OI01
=
3
;
BFMA1O0lOI
=
BFMA1IlI1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:Setup- Burst Mode %0d"
,
BFMA1l01
,
BFMA1O0lOI
)
;
end
5
:
begin
BFMA1OI01
=
3
;
BFMA1I0lOI
=
BFMA1IlI1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:Setup- Alignment %0d"
,
BFMA1l01
,
BFMA1I0lOI
)
;
if
(
BFMA1I0lOI
==
1
|
BFMA1I0lOI
==
2
)
begin
$display
(
"BFM: Untested 8 or 16 Bit alignment selected (WARNING)"
)
;
end
end
6
:
begin
BFMA1OI01
=
3
;
end
7
:
begin
BFMA1OI01
=
3
;
BFMA1l1lOI
=
BFMA1IlI1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:Setup- End Sim Action %0d"
,
BFMA1l01
,
BFMA1l1lOI
)
;
if
(
BFMA1l1lOI
>
2
)
begin
$display
(
"BFM: Unexpected End Simulation value (WARNING)"
)
;
end
end
default
:
begin
$display
(
"BFM Unknown Setup Command (FAILURE)"
)
;
end
endcase
end
BFMA1IOIl
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
BFMA1OI1
<=
(
(
BFMA1lll1
[
1
]
[
0
]
)
==
1
'b
1
)
;
BFMA1II1
<=
(
(
BFMA1lll1
[
1
]
[
1
]
)
==
1
'b
1
)
;
BFMA1lO1
<=
(
(
BFMA1lll1
[
1
]
[
2
]
)
==
1
'b
1
)
;
BFMA1IO1
<=
(
(
BFMA1lll1
[
1
]
[
3
]
)
==
1
'b
1
)
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:drivex %0d "
,
BFMA1l01
,
BFMA1lI
[
1
]
)
;
end
BFMA1IO1I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
3
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:error %0d %0d (No effect in this version)"
,
BFMA1l01
,
BFMA1lI
[
1
]
,
BFMA1lI
[
2
]
)
;
end
BFMA1l10I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
BFMA1I1IOI
=
BFMA1lll1
[
1
]
[
3
:
0
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:prot %0d "
,
BFMA1l01
,
BFMA1I1IOI
)
;
end
BFMA1OO1I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
BFMA1O1IOI
=
BFMA1lll1
[
1
]
[
0
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:lock %0d "
,
BFMA1l01
,
BFMA1O1IOI
)
;
end
BFMA1lO1I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
BFMA1l1IOI
=
BFMA1lll1
[
1
]
[
2
:
0
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:burst %0d "
,
BFMA1l01
,
BFMA1l1IOI
)
;
end
BFMA1OO0I
:
begin
BFMA1OI01
=
2
;
BFMA1lI11
=
BFMA1lI
[
1
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:wait %0d  starting at %0d ns"
,
BFMA1l01
,
BFMA1lI11
,
$time
)
;
BFMA1O001
=
1
;
end
BFMA1OOIl
:
begin
BFMA1OI01
=
2
;
BFMA1O00OI
=
BFMA1lI
[
1
]
*
1000
+
(
$time
/
1
)
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:waitus %0d  starting at %0d ns"
,
BFMA1l01
,
BFMA1lI
[
1
]
,
$time
)
;
BFMA1O001
=
1
;
end
BFMA1l1Ol
:
begin
BFMA1OI01
=
2
;
BFMA1O00OI
=
BFMA1lI
[
1
]
*
1
+
(
$time
/
1
)
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:waitns %0d  starting at %0d ns"
,
BFMA1l01
,
BFMA1lI
[
1
]
,
$time
)
;
BFMA1O001
=
1
;
end
BFMA1OI1I
:
begin
BFMA1OI01
=
3
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:checktime %0d %0d at %0d ns"
,
BFMA1l01
,
BFMA1lI
[
1
]
,
BFMA1lI
[
2
]
,
$time
)
;
BFMA1O001
=
1
;
end
BFMA1lI1I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
1
;
BFMA1l1O1
=
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:starttimer at %0d ns"
,
BFMA1l01
,
$time
)
;
end
BFMA1Ol1I
:
begin
BFMA1OI01
=
3
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:checktimer %0d %0d at %0d ns "
,
BFMA1l01
,
BFMA1lI
[
1
]
,
BFMA1lI
[
2
]
,
$time
)
;
BFMA1O001
=
1
;
end
BFMA1l11
:
begin
BFMA1OI01
=
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:nop"
,
BFMA1l01
)
;
end
BFMA1OOOI
:
begin
BFMA1OI01
=
4
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1Il01
=
BFMA1lll1
[
3
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:write %c %08x %08x at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1Il01
,
$time
)
;
BFMA1I101
=
1
;
end
BFMA1lOII
:
begin
BFMA1OI01
=
5
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1Il01
=
BFMA1lll1
[
3
]
;
BFMA1I00OI
=
BFMA1lll1
[
4
]
[
0
]
;
BFMA1l00OI
=
BFMA1lll1
[
4
]
[
5
:
4
]
;
BFMA1I10OI
=
BFMA1lll1
[
4
]
[
10
:
8
]
;
BFMA1l10OI
=
BFMA1lll1
[
4
]
[
12
]
;
BFMA1O10OI
=
BFMA1lll1
[
4
]
[
19
:
16
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:idle %c %08x %08x %08x at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1Il01
,
BFMA1lll1
[
4
]
,
$time
)
;
BFMA1IO11
=
1
;
end
BFMA1IOOI
:
begin
BFMA1OI01
=
3
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1Il01
=
{
32
{
1
'b
0
}
}
;
BFMA1ll01
=
{
32
{
1
'b
0
}
}
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:read %c %08x at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
$time
)
;
BFMA1I001
=
1
;
end
BFMA1IOII
:
begin
BFMA1OI01
=
4
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1Il01
=
{
32
{
1
'b
0
}
}
;
BFMA1ll01
=
{
32
{
1
'b
0
}
}
;
BFMA1OOlOI
=
BFMA1OOl1
(
BFMA1Ol
[
BFMA1O000
+
3
]
,
BFMA1I01
)
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:readstore %c %08x @%0d at %0d ns "
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1OOlOI
,
$time
)
;
BFMA1I001
=
1
;
BFMA1OO11
=
1
;
end
BFMA1lOOI
:
begin
BFMA1OI01
=
4
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1Il01
=
BFMA1lll1
[
3
]
;
BFMA1ll01
=
{
32
{
1
'b
1
}
}
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:readcheck %c %08x %08x at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1Il01
,
$time
)
;
BFMA1I001
=
1
;
end
BFMA1OIOI
:
begin
BFMA1OI01
=
5
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1Il01
=
BFMA1lll1
[
3
]
;
BFMA1ll01
=
BFMA1lll1
[
4
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:readmask %c %08x %08x %08x at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1Il01
,
BFMA1ll01
,
$time
)
;
BFMA1I001
=
1
;
end
BFMA1IIOI
:
begin
BFMA1OI01
=
4
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1Il01
=
BFMA1lll1
[
3
]
;
BFMA1ll01
=
{
32
{
1
'b
1
}
}
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:poll %c %08x %08x at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1Il01
,
$time
)
;
BFMA1OI11
=
1
;
BFMA1l101
=
1
;
BFMA1l101
=
1
;
end
BFMA1lIOI
:
begin
BFMA1OI01
=
5
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1Il01
=
BFMA1lll1
[
3
]
;
BFMA1ll01
=
BFMA1lll1
[
4
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:pollmask %c %08x %08x %08x at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1Il01
,
BFMA1ll01
,
$time
)
;
BFMA1l101
=
1
;
end
BFMA1OlOI
:
begin
BFMA1OI01
=
5
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1Il01
=
{
32
{
1
'b
0
}
}
;
BFMA1ll01
=
{
32
{
1
'b
0
}
}
;
BFMA1Ol11
=
BFMA1lI
[
3
]
;
BFMA1ll01
[
BFMA1Ol11
]
=
1
'b
1
;
BFMA1Il01
[
BFMA1Ol11
]
=
BFMA1lll1
[
4
]
[
0
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:pollbit %c %08x %0d %0d at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1Ol11
,
BFMA1Il01
[
BFMA1Ol11
]
,
$time
)
;
BFMA1l101
=
1
;
end
BFMA1IlOI
:
begin
BFMA1O111
=
BFMA1lI
[
1
]
;
BFMA1OI01
=
4
+
BFMA1O111
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
2
]
+
BFMA1lI
[
3
]
)
;
BFMA1I111
=
0
;
BFMA1l111
=
BFMA1llO0
(
BFMA1l1l1
,
BFMA1OllOI
)
;
begin
:
BFMA1l11OI
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
BFMA1O111
-
1
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
BFMA1OOOOI
[
BFMA1I0I0
]
=
BFMA1lI
[
BFMA1I0I0
+
4
]
;
end
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:writemultiple %c %08x %08x ... at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1OOOOI
[
0
]
,
$time
)
;
BFMA1l001
=
1
;
end
BFMA1llOI
:
begin
BFMA1O111
=
BFMA1lI
[
3
]
;
BFMA1OI01
=
6
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1I111
=
0
;
BFMA1l111
=
BFMA1llO0
(
BFMA1l1l1
,
BFMA1OllOI
)
;
BFMA1l0OOI
=
BFMA1lI
[
4
]
;
BFMA1O1OOI
=
BFMA1lI
[
5
]
;
begin
:
BFMA1OOOII
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
BFMA1O111
-
1
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
BFMA1OOOOI
[
BFMA1I0I0
]
=
BFMA1l0OOI
;
BFMA1l0OOI
=
BFMA1l0OOI
+
BFMA1O1OOI
;
end
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:fill %c %08x %0d %0d %0d at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1O111
,
BFMA1lI
[
4
]
,
BFMA1lI
[
4
]
,
$time
)
;
BFMA1l001
=
1
;
end
BFMA1O0OI
:
begin
BFMA1O111
=
BFMA1lI
[
4
]
;
BFMA1OI01
=
5
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1I111
=
0
;
BFMA1l111
=
BFMA1llO0
(
BFMA1l1l1
,
BFMA1OllOI
)
;
BFMA1lIOOI
=
BFMA1lI
[
3
]
;
begin
:
BFMA1IOOII
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
BFMA1O111
-
1
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
BFMA1OOOOI
[
BFMA1I0I0
]
=
BFMA1Ol
[
2
+
BFMA1lIOOI
+
BFMA1I0I0
]
;
end
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:writetable %c %08x %0d %0d at %0d ns "
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1lIOOI
,
BFMA1O111
,
$time
)
;
BFMA1l001
=
1
;
end
BFMA1OIII
:
begin
BFMA1O111
=
BFMA1lI
[
4
]
;
BFMA1OI01
=
5
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1I111
=
0
;
BFMA1l111
=
BFMA1llO0
(
BFMA1l1l1
,
BFMA1OllOI
)
;
BFMA1lOIOI
=
BFMA1OOl1
(
BFMA1Ol
[
BFMA1O000
+
3
]
,
BFMA1I01
)
;
begin
:
BFMA1lOOII
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
BFMA1O111
-
1
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
BFMA1OOOOI
[
BFMA1I0I0
]
=
BFMA1ll1
[
BFMA1lOIOI
+
BFMA1I0I0
]
;
end
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:writearray %c %08x %0d %0d at %0d ns "
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1lOIOI
,
BFMA1O111
,
$time
)
;
BFMA1l001
=
1
;
end
BFMA1I0OI
:
begin
BFMA1O111
=
BFMA1lI
[
3
]
;
BFMA1OI01
=
4
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1ll01
=
{
32
{
1
'b
0
}
}
;
BFMA1I111
=
0
;
BFMA1l111
=
BFMA1llO0
(
BFMA1l1l1
,
BFMA1OllOI
)
;
BFMA1ll01
=
{
32
{
1
'b
0
}
}
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:readmult %c %08x %0d at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1O111
,
$time
)
;
BFMA1O101
=
1
;
end
BFMA1l0OI
:
begin
BFMA1O111
=
BFMA1lI
[
1
]
;
BFMA1OI01
=
4
+
BFMA1O111
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
2
]
+
BFMA1lI
[
3
]
)
;
BFMA1ll01
=
{
32
{
1
'b
1
}
}
;
BFMA1I111
=
0
;
BFMA1l111
=
BFMA1llO0
(
BFMA1l1l1
,
BFMA1OllOI
)
;
BFMA1ll01
=
{
32
{
1
'b
1
}
}
;
begin
:
BFMA1OIOII
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
BFMA1O111
-
1
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
BFMA1OOOOI
[
BFMA1I0I0
]
=
BFMA1lI
[
BFMA1I0I0
+
4
]
;
end
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:readmultchk %c %08x %08x ... at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1OOOOI
[
0
]
,
$time
)
;
BFMA1O101
=
1
;
end
BFMA1O1OI
:
begin
BFMA1O111
=
BFMA1lI
[
3
]
;
BFMA1OI01
=
6
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1ll01
=
{
32
{
1
'b
1
}
}
;
BFMA1I111
=
0
;
BFMA1l111
=
BFMA1llO0
(
BFMA1l1l1
,
BFMA1OllOI
)
;
BFMA1l0OOI
=
BFMA1lI
[
4
]
;
BFMA1O1OOI
=
BFMA1lI
[
5
]
;
begin
:
BFMA1IIOII
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
BFMA1O111
-
1
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
BFMA1OOOOI
[
BFMA1I0I0
]
=
BFMA1l0OOI
;
BFMA1l0OOI
=
BFMA1l0OOI
+
BFMA1O1OOI
;
end
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:fillcheck %c %08x %0d %0d %0d at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1O111
,
BFMA1lI
[
4
]
,
BFMA1lI
[
5
]
,
$time
)
;
BFMA1O101
=
1
;
end
BFMA1I1OI
:
begin
BFMA1O111
=
BFMA1lI
[
4
]
;
BFMA1OI01
=
5
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1ll01
=
{
32
{
1
'b
1
}
}
;
BFMA1I111
=
0
;
BFMA1l111
=
BFMA1llO0
(
BFMA1l1l1
,
BFMA1OllOI
)
;
BFMA1lIOOI
=
BFMA1lI
[
3
]
;
begin
:
BFMA1lIOII
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
BFMA1O111
-
1
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
BFMA1OOOOI
[
BFMA1I0I0
]
=
BFMA1Ol
[
BFMA1lIOOI
+
2
+
BFMA1I0I0
]
;
end
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:readtable %c %08x %0d %0d at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1lIOOI
,
BFMA1O111
,
$time
)
;
BFMA1O101
=
1
;
end
BFMA1IIII
:
begin
BFMA1O111
=
BFMA1lI
[
4
]
;
BFMA1OI01
=
5
;
BFMA1lI01
=
BFMA1I0O0
(
BFMA1l1l1
,
BFMA1lIlOI
)
;
BFMA1Ol01
=
to_slv32
(
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
)
;
BFMA1ll01
=
{
32
{
1
'b
1
}
}
;
BFMA1I111
=
0
;
BFMA1l111
=
BFMA1llO0
(
BFMA1l1l1
,
BFMA1OllOI
)
;
BFMA1lOIOI
=
BFMA1OOl1
(
BFMA1Ol
[
BFMA1O000
+
3
]
,
BFMA1I01
)
;
begin
:
BFMA1OlOII
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
BFMA1O111
-
1
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
BFMA1OOOOI
[
BFMA1I0I0
]
=
BFMA1ll1
[
BFMA1lOIOI
+
BFMA1I0I0
]
;
end
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:readtable %c %08x %0d %0d at %0d ns"
,
BFMA1l01
,
BFMA1IlO0
(
BFMA1l1l1
)
,
BFMA1Ol01
,
BFMA1lOIOI
,
BFMA1O111
,
$time
)
;
BFMA1O101
=
1
;
end
BFMA1O00I
:
begin
BFMA1OI01
=
7
;
BFMA1O001
=
1
;
BFMA1lOO1
=
BFMA1Il10
;
end
BFMA1I00I
:
begin
BFMA1OI01
=
7
;
BFMA1O001
=
1
;
BFMA1lOO1
=
BFMA1Il10
;
end
BFMA1O1II
:
begin
BFMA1OI01
=
1
;
BFMA1IlOOI
=
0
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:waitfiq at %0d ns "
,
BFMA1l01
,
$time
)
;
BFMA1O001
=
1
;
end
BFMA1I1II
:
begin
BFMA1OI01
=
1
;
BFMA1IlOOI
=
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:waitirq at %0d ns "
,
BFMA1l01
,
$time
)
;
BFMA1O001
=
1
;
end
BFMA1l0II
:
begin
BFMA1OI01
=
2
;
BFMA1IlOOI
=
BFMA1lI
[
1
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:waitint %0d  at %0d ns"
,
BFMA1l01
,
BFMA1IlOOI
,
$time
)
;
BFMA1O001
=
1
;
end
BFMA1lIII
:
begin
BFMA1OI01
=
2
;
BFMA1Il01
=
BFMA1lll1
[
1
]
;
BFMA1O10
<=
BFMA1Il01
;
BFMA1OO0
<=
1
'b
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:iowrite %08x  at %0d ns "
,
BFMA1l01
,
BFMA1Il01
,
$time
)
;
end
BFMA1OlII
:
begin
BFMA1OI01
=
2
;
BFMA1Il01
=
{
32
{
1
'b
0
}
}
;
BFMA1ll01
=
{
32
{
1
'b
0
}
}
;
BFMA1OOlOI
=
BFMA1OOl1
(
BFMA1Ol
[
BFMA1O000
+
1
]
,
BFMA1I01
)
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:ioread @%0d at %0d ns"
,
BFMA1l01
,
BFMA1OOlOI
,
$time
)
;
BFMA1l1l
<=
1
'b
1
;
BFMA1O001
=
1
;
BFMA1OO11
=
1
;
BFMA1lO11
=
1
;
end
BFMA1IlII
:
begin
BFMA1OI01
=
2
;
BFMA1Il01
=
BFMA1lll1
[
1
]
;
BFMA1ll01
=
{
32
{
1
'b
1
}
}
;
BFMA1l1l
<=
1
'b
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:iocheck %08x  at %0d ns "
,
BFMA1l01
,
BFMA1Il01
,
$time
)
;
BFMA1O001
=
1
;
end
BFMA1llII
:
begin
BFMA1OI01
=
3
;
BFMA1Il01
=
BFMA1lll1
[
1
]
;
BFMA1ll01
=
BFMA1lll1
[
2
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:iomask %08x %08x  at %0d ns"
,
BFMA1l01
,
BFMA1Il01
,
BFMA1ll01
,
$time
)
;
BFMA1l1l
<=
1
'b
1
;
BFMA1O001
=
1
;
end
BFMA1l1OI
:
begin
BFMA1OI01
=
2
;
BFMA1Il01
=
{
32
{
1
'b
0
}
}
;
BFMA1ll01
=
{
32
{
1
'b
0
}
}
;
BFMA1Ol11
=
BFMA1lI
[
1
]
;
BFMA1Il01
[
BFMA1Ol11
]
=
BFMA1I1l1
[
0
]
;
BFMA1ll01
[
BFMA1Ol11
]
=
1
'b
1
;
BFMA1l1l
<=
1
'b
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:iotest %0d %0d  at %0d ns"
,
BFMA1l01
,
BFMA1Ol11
,
BFMA1I1l1
[
0
]
,
$time
)
;
BFMA1O001
=
1
;
end
BFMA1O0II
:
begin
BFMA1OI01
=
2
;
BFMA1Ol11
=
BFMA1lI
[
1
]
;
BFMA1O10
[
BFMA1Ol11
]
<=
1
'b
1
;
BFMA1OO0
<=
1
'b
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:ioset %0d at %0d ns"
,
BFMA1l01
,
BFMA1Ol11
,
$time
)
;
end
BFMA1I0II
:
begin
BFMA1OI01
=
2
;
BFMA1Ol11
=
BFMA1lI
[
1
]
;
BFMA1O10
[
BFMA1Ol11
]
<=
1
'b
0
;
BFMA1OO0
<=
1
'b
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:ioclr %0d at %0d ns"
,
BFMA1l01
,
BFMA1Ol11
,
$time
)
;
end
BFMA1OOII
:
begin
BFMA1OI01
=
2
;
BFMA1Il01
=
{
32
{
1
'b
0
}
}
;
BFMA1ll01
=
{
32
{
1
'b
0
}
}
;
BFMA1Ol11
=
BFMA1lI
[
1
]
;
BFMA1Il01
[
BFMA1Ol11
]
=
BFMA1I1l1
[
0
]
;
BFMA1ll01
[
BFMA1Ol11
]
=
1
'b
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:iowait %0d %0d at %0d ns "
,
BFMA1l01
,
BFMA1Ol11
,
BFMA1I1l1
[
0
]
,
$time
)
;
BFMA1l1l
<=
1
'b
1
;
BFMA1O001
=
1
;
end
BFMA1OOlI
:
begin
BFMA1OI01
=
3
;
BFMA1Ol01
=
BFMA1lll1
[
1
]
;
BFMA1Il01
=
BFMA1lll1
[
2
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:extwrite %08x %08x at %0d ns"
,
BFMA1l01
,
BFMA1Ol01
,
BFMA1Il01
,
$time
)
;
BFMA1O001
=
1
;
end
BFMA1IOlI
:
begin
BFMA1OI01
=
3
;
BFMA1Ol01
=
BFMA1lll1
[
1
]
;
BFMA1Il01
=
{
32
{
1
'b
0
}
}
;
BFMA1ll01
=
{
32
{
1
'b
0
}
}
;
BFMA1OOlOI
=
BFMA1OOl1
(
BFMA1Ol
[
BFMA1O000
+
2
]
,
BFMA1I01
)
;
BFMA1O1l
<=
1
'b
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:extread @%0d %08x at %0d ns "
,
BFMA1l01
,
BFMA1OOlOI
,
BFMA1Ol01
,
$time
)
;
BFMA1O001
=
1
;
BFMA1OO11
=
1
;
BFMA1lO11
=
1
;
end
BFMA1lIlI
:
begin
BFMA1O111
=
BFMA1lI
[
1
]
;
BFMA1l011
=
BFMA1lI
[
2
]
;
BFMA1OI01
=
BFMA1O111
+
3
;
begin
:
BFMA1IlOII
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<
BFMA1O111
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
BFMA1OOOOI
[
BFMA1I0I0
]
=
BFMA1lI
[
BFMA1I0I0
+
3
]
;
end
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:extwrite %08x %0d Words at %0t ns"
,
BFMA1l01
,
BFMA1Ol01
,
BFMA1O111
,
$time
)
;
BFMA1I111
=
0
;
BFMA1O001
=
1
;
end
BFMA1lOlI
:
begin
BFMA1OI01
=
3
;
BFMA1Ol01
=
BFMA1lll1
[
1
]
;
BFMA1Il01
=
BFMA1lll1
[
2
]
;
BFMA1ll01
=
{
32
{
1
'b
1
}
}
;
BFMA1OI11
=
1
;
BFMA1O1l
<=
1
'b
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:extcheck %08x %08x at %0d ns"
,
BFMA1l01
,
BFMA1Ol01
,
BFMA1Il01
,
$time
)
;
BFMA1O001
=
1
;
end
BFMA1OIlI
:
begin
BFMA1OI01
=
4
;
BFMA1Ol01
=
BFMA1lll1
[
1
]
;
BFMA1Il01
=
BFMA1lll1
[
2
]
;
BFMA1ll01
=
BFMA1lll1
[
3
]
;
BFMA1O1l
<=
1
'b
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:extmask %08x %08x %08x at %0d ns"
,
BFMA1l01
,
BFMA1Ol01
,
BFMA1Il01
,
BFMA1ll01
,
$time
)
;
BFMA1O001
=
1
;
end
BFMA1IIlI
:
begin
BFMA1OI01
=
1
;
BFMA1lI11
=
1
;
BFMA1OI11
=
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:extwait "
,
BFMA1l01
)
;
BFMA1O001
=
1
;
end
BFMA1OllI
:
begin
$display
(
"LABEL instructions not allowed in vector files (FAILURE)"
)
;
end
BFMA1II0I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
+
BFMA1lI
[
1
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:table %08x ... (length=%0d)"
,
BFMA1l01
,
BFMA1lI
[
2
]
,
BFMA1OI01
-
2
)
;
end
BFMA1IllI
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
BFMA1I0OOI
=
BFMA1lI
[
1
]
;
BFMA1OI01
=
BFMA1I0OOI
-
BFMA1O000
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:jump"
,
BFMA1l01
)
;
end
BFMA1lllI
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
3
;
BFMA1I0OOI
=
BFMA1lI
[
1
]
;
if
(
BFMA1lI
[
2
]
==
0
)
begin
BFMA1OI01
=
BFMA1I0OOI
-
BFMA1O000
;
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:jumpz  %08x"
,
BFMA1l01
,
BFMA1lI
[
2
]
)
;
end
BFMA1lOOl
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
5
;
BFMA1I0OOI
=
BFMA1lI
[
1
]
;
BFMA1OIIOI
=
BFMA1O1O0
(
BFMA1lI
[
3
]
,
BFMA1lI
[
2
]
,
BFMA1lI
[
4
]
,
DEBUG
)
;
if
(
BFMA1OIIOI
==
0
)
begin
BFMA1OI01
=
BFMA1I0OOI
+
2
-
BFMA1O000
;
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:if %08x func %08x"
,
BFMA1l01
,
BFMA1lI
[
2
]
,
BFMA1lI
[
4
]
)
;
end
BFMA1OIOl
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
5
;
BFMA1I0OOI
=
BFMA1lI
[
1
]
;
BFMA1OIIOI
=
BFMA1O1O0
(
BFMA1lI
[
3
]
,
BFMA1lI
[
2
]
,
BFMA1lI
[
4
]
,
DEBUG
)
;
if
(
BFMA1OIIOI
!=
0
)
begin
BFMA1OI01
=
BFMA1I0OOI
+
2
-
BFMA1O000
;
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:ifnot %08x func %08x"
,
BFMA1l01
,
BFMA1lI
[
2
]
,
BFMA1lI
[
4
]
)
;
end
BFMA1lIOl
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
BFMA1I0OOI
=
BFMA1lI
[
1
]
;
BFMA1OI01
=
BFMA1I0OOI
+
2
-
BFMA1O000
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:else "
,
BFMA1l01
)
;
end
BFMA1OlOl
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:endif "
,
BFMA1l01
)
;
end
BFMA1IIOl
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
5
;
BFMA1I0OOI
=
BFMA1lI
[
1
]
+
2
;
BFMA1OIIOI
=
BFMA1O1O0
(
BFMA1lI
[
3
]
,
BFMA1lI
[
2
]
,
BFMA1lI
[
4
]
,
DEBUG
)
;
if
(
BFMA1OIIOI
==
0
)
begin
BFMA1OI01
=
BFMA1I0OOI
-
BFMA1O000
;
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:while %08x func %08x"
,
BFMA1l01
,
BFMA1lI
[
2
]
,
BFMA1lI
[
4
]
)
;
end
BFMA1IlOl
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
BFMA1I0OOI
=
BFMA1lI
[
1
]
;
BFMA1OI01
=
BFMA1I0OOI
-
BFMA1O000
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:endwhile"
,
BFMA1l01
)
;
end
BFMA1O0Ol
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
4
;
BFMA1I0OOI
=
BFMA1lI
[
3
]
;
if
(
BFMA1lI
[
1
]
!=
BFMA1lI
[
2
]
)
begin
BFMA1OI01
=
BFMA1I0OOI
-
BFMA1O000
;
end
else
begin
BFMA1O01OI
[
BFMA1I01OI
]
=
1
;
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:when %08x=%08x %08x"
,
BFMA1l01
,
BFMA1lI
[
1
]
,
BFMA1lI
[
2
]
,
BFMA1lI
[
3
]
)
;
end
BFMA1l0Ol
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
4
;
BFMA1I0OOI
=
BFMA1lI
[
3
]
;
if
(
BFMA1O01OI
[
BFMA1I01OI
]
)
begin
BFMA1OI01
=
BFMA1I0OOI
-
BFMA1O000
;
end
else
begin
BFMA1O01OI
[
BFMA1I01OI
]
=
0
;
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:default %08x=%08x %08x"
,
BFMA1l01
,
BFMA1lI
[
1
]
,
BFMA1lI
[
2
]
,
BFMA1lI
[
3
]
)
;
end
BFMA1llOl
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
1
;
BFMA1I01OI
=
BFMA1I01OI
+
1
;
BFMA1O01OI
[
BFMA1I01OI
]
=
0
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:case"
,
BFMA1l01
)
;
end
BFMA1I0Ol
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
1
;
BFMA1I01OI
=
BFMA1I01OI
-
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:endcase"
,
BFMA1l01
)
;
end
BFMA1O0lI
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
3
;
BFMA1I0OOI
=
BFMA1lI
[
1
]
;
if
(
BFMA1lI
[
2
]
!=
0
)
begin
BFMA1OI01
=
BFMA1I0OOI
-
BFMA1O000
;
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:jumpnz  %08x"
,
BFMA1l01
,
BFMA1lI
[
2
]
)
;
end
BFMA1l11I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
4
;
BFMA1Il01
=
BFMA1lll1
[
2
]
;
BFMA1ll01
=
BFMA1lll1
[
3
]
;
BFMA1Il0OI
=
(
BFMA1lll1
[
1
]
^
BFMA1Il01
)
&
BFMA1ll01
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:compare  %08x==%08x Mask=%08x (RES=%08x) at %0d ns"
,
BFMA1l01
,
BFMA1lI
[
1
]
,
BFMA1Il01
,
BFMA1ll01
,
BFMA1Il0OI
,
$time
)
;
if
(
BFMA1Il0OI
!=
0
)
begin
BFMA1II10
=
BFMA1II10
+
1
;
$display
(
"ERROR:  compare failed %08x==%08x Mask=%08x (RES=%08x) "
,
BFMA1lI
[
1
]
,
BFMA1Il01
,
BFMA1ll01
,
BFMA1Il0OI
)
;
$display
(
"       Stimulus file %0s  Line No %0d"
,
BFMA1lOlOI
[
BFMA1OIl0
(
BFMA1l01
,
BFMA1IIlOI
)
]
,
BFMA1l1I0
(
BFMA1l01
,
BFMA1IIlOI
)
)
;
$display
(
"BFM Data Compare Error (ERROR)"
)
;
$stop
;
end
end
BFMA1O1Ol
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
4
;
BFMA1Il01
=
BFMA1lll1
[
2
]
;
BFMA1ll01
=
BFMA1lll1
[
3
]
;
if
(
BFMA1lI
[
1
]
>=
BFMA1lI
[
2
]
&
BFMA1lI
[
1
]
<=
BFMA1lI
[
3
]
)
begin
BFMA1Il0OI
=
1
;
end
else
begin
BFMA1Il0OI
=
0
;
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:cmprange %0d in %0d to %0d at %0d ns"
,
BFMA1l01
,
BFMA1lI
[
1
]
,
BFMA1lI
[
2
]
,
BFMA1lI
[
3
]
,
$time
)
;
if
(
BFMA1Il0OI
==
0
)
begin
BFMA1II10
=
BFMA1II10
+
1
;
$display
(
"ERROR: cmprange failed %0d in %0d to %0d"
,
BFMA1lI
[
1
]
,
BFMA1lI
[
2
]
,
BFMA1lI
[
3
]
)
;
$display
(
"       Stimulus file %0s  Line No %0d"
,
BFMA1lOlOI
[
BFMA1OIl0
(
BFMA1l01
,
BFMA1IIlOI
)
]
,
BFMA1l1I0
(
BFMA1l01
,
BFMA1IIlOI
)
)
;
$display
(
"BFM Data Compare Error (ERROR)"
)
;
$stop
;
end
end
BFMA1O11I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
BFMA1lI00
=
BFMA1lI
[
1
]
;
BFMA1I01
=
BFMA1I01
+
BFMA1lI00
;
BFMA1ll1
[
BFMA1I01
]
=
0
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:int %0d"
,
BFMA1l01
,
BFMA1lI
[
1
]
)
;
end
BFMA1I0lI
,
BFMA1l0lI
:
begin
BFMA1OI1OI
=
1
;
if
(
BFMA1OO01
==
BFMA1I0lI
)
begin
BFMA1OI01
=
2
;
BFMA1lI00
=
0
;
end
else
begin
BFMA1lI00
=
BFMA1lI
[
2
]
;
BFMA1OI01
=
3
+
BFMA1lI00
;
end
BFMA1llOOI
=
BFMA1lI
[
1
]
;
BFMA1O0OOI
=
BFMA1O000
+
BFMA1OI01
;
BFMA1OI01
=
BFMA1llOOI
-
BFMA1O000
;
BFMA1ll1
[
BFMA1I01
]
=
BFMA1O0OOI
;
BFMA1I01
=
BFMA1I01
+
1
;
if
(
BFMA1lI00
>
0
)
begin
begin
:
BFMA1llOII
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
BFMA1lI00
-
1
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
BFMA1ll1
[
BFMA1I01
]
=
BFMA1lI
[
3
+
BFMA1I0I0
]
;
BFMA1I01
=
BFMA1I01
+
1
;
end
end
end
if
(
DEBUG
>=
2
&
BFMA1OO01
==
BFMA1I0lI
)
$display
(
"BFM:%0d:call %0d"
,
BFMA1l01
,
BFMA1llOOI
)
;
if
(
DEBUG
>=
2
&
BFMA1OO01
==
BFMA1l0lI
)
$display
(
"BFM:%0d:call %0d %08x ..."
,
BFMA1l01
,
BFMA1llOOI
,
BFMA1lI
[
3
]
)
;
end
BFMA1O1lI
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
BFMA1I01
=
BFMA1I01
-
BFMA1lI
[
1
]
;
BFMA1O0OOI
=
0
;
if
(
BFMA1I01
>
0
)
begin
BFMA1I01
=
BFMA1I01
-
1
;
BFMA1O0OOI
=
BFMA1ll1
[
BFMA1I01
]
;
end
if
(
BFMA1O0OOI
==
0
)
begin
BFMA1lOOOI
=
1
;
BFMA1OO11
=
1
;
BFMA1OI1OI
=
0
;
end
else
begin
BFMA1OI01
=
BFMA1O0OOI
-
BFMA1O000
;
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:return"
,
BFMA1l01
)
;
end
BFMA1I1Ol
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
3
;
BFMA1I01
=
BFMA1I01
-
BFMA1lI
[
1
]
;
BFMA1O0OOI
=
0
;
if
(
BFMA1I01
>
0
)
begin
BFMA1I01
=
BFMA1I01
-
1
;
BFMA1O0OOI
=
BFMA1ll1
[
BFMA1I01
]
;
end
BFMA1O01
=
BFMA1lI
[
2
]
;
if
(
BFMA1O0OOI
==
0
)
begin
BFMA1lOOOI
=
1
;
BFMA1OO11
=
1
;
BFMA1OI1OI
=
0
;
end
else
begin
BFMA1OI01
=
BFMA1O0OOI
-
BFMA1O000
;
end
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:return %08x"
,
BFMA1l01
,
BFMA1O01
)
;
end
BFMA1I1lI
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
5
;
BFMA1lOIOI
=
BFMA1OOl1
(
BFMA1Ol
[
BFMA1O000
+
1
]
,
BFMA1I01
)
;
BFMA1OIIOI
=
BFMA1lI
[
2
]
;
BFMA1ll1
[
BFMA1lOIOI
]
=
BFMA1OIIOI
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:loop %0d %0d %0d %0d "
,
BFMA1l01
,
BFMA1lOIOI
,
BFMA1lI
[
2
]
,
BFMA1lI
[
3
]
,
BFMA1lI
[
4
]
)
;
end
BFMA1l1lI
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
BFMA1I0l1
=
BFMA1lI
[
1
]
;
begin
:
BFMA1O0OII
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
2
;
BFMA1I0I0
<=
4
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
BFMA1Ill1
[
BFMA1I0I0
]
=
BFMA1lII1
(
(
to_slv32
(
BFMA1Ol
[
BFMA1I0l1
]
[
7
+
BFMA1I0I0
]
)
==
1
'b
1
)
,
BFMA1Ol
[
BFMA1I0l1
+
BFMA1I0I0
]
)
;
end
end
BFMA1lOIOI
=
BFMA1OOl1
(
BFMA1Ol
[
BFMA1I0l1
+
1
]
,
BFMA1I01
)
;
BFMA1Il00
=
BFMA1Ill1
[
4
]
;
BFMA1I100
=
BFMA1Ill1
[
3
]
;
BFMA1O1l1
=
BFMA1ll1
[
BFMA1lOIOI
]
;
BFMA1O1l1
=
BFMA1O1l1
+
BFMA1Il00
;
BFMA1ll1
[
BFMA1lOIOI
]
=
BFMA1O1l1
;
BFMA1I0OOI
=
BFMA1I0l1
+
5
;
if
(
(
BFMA1Il00
>=
0
&
BFMA1O1l1
<=
BFMA1I100
)
|
(
BFMA1Il00
<
0
&
BFMA1O1l1
>=
BFMA1I100
)
)
begin
BFMA1OI01
=
BFMA1I0OOI
-
BFMA1O000
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:endloop (Next Loop=%0d)"
,
BFMA1l01
,
BFMA1O1l1
)
;
end
else
begin
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:endloop (Finished)"
,
BFMA1l01
)
;
end
end
BFMA1OI0I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
BFMA1II01
=
BFMA1lI
[
1
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:timeout %0d"
,
BFMA1l01
,
BFMA1II01
)
;
end
BFMA1Il1I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
BFMA1lO10
=
BFMA1lI
[
1
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:rand %0d"
,
BFMA1l01
,
BFMA1lO10
)
;
end
BFMA1Ol0I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
BFMA1OI00
(
BFMA1Ol
[
BFMA1O000
+
1
]
)
;
BFMA1l000
=
BFMA1ll00
(
BFMA1O000
)
;
$display
(
"BFM:%0s"
,
BFMA1l000
)
;
end
BFMA1Il0I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
BFMA1OI00
(
BFMA1Ol
[
BFMA1O000
+
1
]
)
;
BFMA1l000
=
BFMA1ll00
(
BFMA1O000
)
;
$display
(
"################################################################"
)
;
$display
(
"BFM:%0s"
,
BFMA1l000
)
;
end
BFMA1ll0I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OlOOI
=
BFMA1O01l
(
BFMA1I1l1
[
15
:
8
]
)
;
BFMA1OI01
=
(
BFMA1OlOOI
-
1
)
/
4
+
2
;
end
BFMA1I10I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
if
(
DEBUGLEVEL
>=
0
&
DEBUGLEVEL
<=
5
)
begin
$display
(
"BFM:%0d: DEBUG - ignored due to DEBUGLEVEL generic setting"
,
BFMA1l01
)
;
end
else
begin
DEBUG
<=
BFMA1lI
[
1
]
;
$display
(
"BFM:%0d: DEBUG %0d"
,
BFMA1l01
,
BFMA1lI
[
1
]
)
;
end
end
BFMA1l1II
:
begin
BFMA1OI1OI
=
0
;
BFMA1OI01
=
2
;
BFMA1I1OOI
=
BFMA1lI
[
1
]
;
BFMA1l0IOI
[
1
]
=
BFMA1OI
;
if
(
BFMA1I1OOI
==
2
)
begin
if
(
BFMA1O0IOI
)
begin
BFMA1l0IOI
[
1
:
9
]
=
{
"OCCURRED"
,
BFMA1OI
}
;
end
else
begin
$display
(
"BFM: HRESP Did Not Occur When Expected (ERROR)"
)
;
BFMA1II10
=
BFMA1II10
+
1
;
$stop
;
end
BFMA1I1OOI
=
0
;
end
BFMA1O0IOI
=
0
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:hresp %0d %0s"
,
BFMA1l01
,
BFMA1I1OOI
,
BFMA1l0IOI
)
;
end
BFMA1IO0I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:stop %0d"
,
BFMA1l01
,
BFMA1lI
[
1
]
)
;
$display
(
"       Stimulus file %0s  Line No %0d"
,
BFMA1lOlOI
[
BFMA1OIl0
(
BFMA1l01
,
BFMA1IIlOI
)
]
,
BFMA1l1I0
(
BFMA1l01
,
BFMA1IIlOI
)
)
;
case
(
BFMA1lI
[
1
]
)
0
:
begin
$display
(
"BFM Script Stop Command (NOTE)"
)
;
end
1
:
begin
$display
(
"BFM Script Stop Command (WARNING)"
)
;
end
3
:
begin
$display
(
"BFM Script Stop Command (FAILURE)"
)
;
$stop
;
end
default
:
begin
$display
(
"BFM Script Stop Command (ERROR)"
)
;
$stop
;
end
endcase
end
BFMA1lO0I
:
begin
BFMA1lOOOI
=
1
;
end
BFMA1OlIl
:
begin
BFMA1OI1OI
=
1
;
if
(
DEBUG
>=
1
)
$display
(
"BFM:%0d:echo at %0d ns"
,
BFMA1l01
,
$time
)
;
BFMA1OI01
=
2
+
BFMA1lI
[
1
]
;
$display
(
"BFM Parameter values are"
)
;
begin
:
BFMA1I0OII
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
BFMA1OI01
-
3
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
$display
(
" Para %0d=0x%08x (%0d)"
,
BFMA1I0I0
+
1
,
BFMA1lll1
[
2
+
BFMA1I0I0
]
,
BFMA1lll1
[
2
+
BFMA1I0I0
]
)
;
end
end
end
BFMA1lI0I
:
begin
BFMA1OI01
=
2
;
BFMA1lI11
=
BFMA1lI
[
1
]
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:flush %0d at %0d ns"
,
BFMA1l01
,
BFMA1lI11
,
$time
)
;
BFMA1OO11
=
1
;
BFMA1O001
=
1
;
end
BFMA1II1I
:
begin
BFMA1OI1OI
=
1
;
BFMA1II10
=
BFMA1II10
+
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:setfail"
,
BFMA1l01
)
;
$display
(
"BFM: User Script detected ERROR (ERROR)"
)
;
$stop
;
end
BFMA1I01I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
3
;
BFMA1lOIOI
=
BFMA1OOl1
(
BFMA1Ol
[
BFMA1O000
+
1
]
,
BFMA1I01
)
;
BFMA1OIIOI
=
BFMA1lI
[
2
]
;
BFMA1ll1
[
BFMA1lOIOI
]
=
BFMA1OIIOI
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:set %0d= 0x%08x (%0d)"
,
BFMA1l01
,
BFMA1lOIOI
,
BFMA1OIIOI
,
BFMA1OIIOI
)
;
end
BFMA1I11I
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
BFMA1lI
[
2
]
+
3
;
BFMA1lOIOI
=
BFMA1OOl1
(
BFMA1Ol
[
BFMA1O000
+
1
]
,
BFMA1I01
)
;
BFMA1OIIOI
=
BFMA1O1O0
(
BFMA1lI
[
4
]
,
BFMA1lI
[
3
]
,
BFMA1lI
[
5
]
,
DEBUG
)
;
BFMA1I0I0
=
6
;
while
(
BFMA1I0I0
<
BFMA1OI01
)
begin
BFMA1OIIOI
=
BFMA1O1O0
(
BFMA1lI
[
BFMA1I0I0
]
,
BFMA1OIIOI
,
BFMA1lI
[
BFMA1I0I0
+
1
]
,
DEBUG
)
;
BFMA1I0I0
=
BFMA1I0I0
+
2
;
end
BFMA1ll1
[
BFMA1lOIOI
]
=
BFMA1OIIOI
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:set %0d= 0x%08x (%0d)"
,
BFMA1l01
,
BFMA1lOIOI
,
BFMA1OIIOI
,
BFMA1OIIOI
)
;
end
BFMA1OIIl
:
begin
BFMA1OI1OI
=
1
;
if
(
BFMA1O11
)
begin
$fflush
(
BFMA1lIl1
)
;
$fclose
(
BFMA1lIl1
)
;
end
BFMA1OI01
=
BFMA1OI00
(
BFMA1Ol
[
BFMA1O000
+
1
]
)
;
BFMA1I011
=
BFMA1ll00
(
BFMA1O000
)
;
$display
(
"BFM:%0d:LOGFILE %0s"
,
BFMA1l01
,
BFMA1I011
)
;
BFMA1lIl1
=
$fopen
(
BFMA1I011
,
"w"
)
;
BFMA1O11
=
1
;
end
BFMA1IIIl
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
2
;
$display
(
"BFM:%0d:LOGSTART %0d"
,
BFMA1l01
,
BFMA1lI
[
1
]
)
;
if
(
BFMA1O11
==
0
)
begin
$display
(
"Logfile not defined, ignoring command (ERROR)"
)
;
end
else
begin
BFMA1lO0OI
=
(
(
BFMA1lll1
[
1
]
[
0
]
)
==
1
'b
1
)
;
BFMA1OI0OI
=
(
(
BFMA1lll1
[
1
]
[
1
]
)
==
1
'b
1
)
;
BFMA1II0OI
=
(
(
BFMA1lll1
[
1
]
[
2
]
)
==
1
'b
1
)
;
BFMA1lI0OI
=
(
(
BFMA1lll1
[
1
]
[
3
]
)
==
1
'b
1
)
;
end
end
BFMA1lIIl
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
1
;
$display
(
"BFM:%0d:LOGSTOP"
,
BFMA1l01
)
;
BFMA1lO0OI
=
0
;
BFMA1OI0OI
=
0
;
BFMA1II0OI
=
0
;
BFMA1lI0OI
=
0
;
end
BFMA1lOIl
:
begin
BFMA1OI1OI
=
1
;
BFMA1OI01
=
1
;
$display
(
"BFM:%0d:VERSION"
,
BFMA1l01
)
;
$display
(
"  BFM Verilog Version %0s"
,
BFMA1O
)
;
$display
(
"  BFM Date %0s"
,
BFMA1I
)
;
$display
(
"  SVN Revision $Revision: 6419 $"
)
;
$display
(
"  SVN Date $Date: 2009-02-04 04:34:22 -0800 (Wed, 04 Feb 2009) $"
)
;
$display
(
"  Compiler Version %0d"
,
BFMA1Ol0OI
)
;
$display
(
"  Vectors Version %0d"
,
BFMA1ll0OI
)
;
$display
(
"  No of Vectors %0d"
,
BFMA1O0l1
)
;
if
(
BFMA1O11
!=
BFMA1OI
)
begin
$fdisplay
(
BFMA1lIl1
,
"%05d VR %0s %0s %0d %0d %0d"
,
$time
,
BFMA1O
,
BFMA1I
,
BFMA1Ol0OI
,
BFMA1ll0OI
,
BFMA1O0l1
)
;
end
end
default
:
begin
$display
(
"BFM: Instruction %0d Line Number %0d Command %0d"
,
BFMA1O000
,
BFMA1l01
,
BFMA1OO01
)
;
$display
(
"       Stimulus file %0s  Line No %0d"
,
BFMA1lOlOI
[
BFMA1OIl0
(
BFMA1l01
,
BFMA1IIlOI
)
]
,
BFMA1l1I0
(
BFMA1l01
,
BFMA1IIlOI
)
)
;
$display
(
"Instruction not yet implemented (ERROR)"
)
;
$stop
;
end
endcase
end
if
(
BFMA1OI1OI
)
begin
BFMA1OI11
=
0
;
BFMA1O000
=
BFMA1O000
+
BFMA1OI01
;
BFMA1OI01
=
0
;
end
end
BFMA1OlIOI
=
0
;
BFMA1IlIOI
=
0
;
BFMA1llIOI
=
0
;
if
(
BFMA1IlI
==
1
'b
1
)
begin
BFMA1IIIOI
=
BFMA1OOl
&
BFMA1IOl
;
BFMA1lIIOI
=
HRDATA
&
BFMA1IOl
;
BFMA1OlIOI
=
(
BFMA1IIIOI
===
BFMA1lIIOI
)
;
end
if
(
BFMA1I1l
==
1
'b
1
)
begin
BFMA1IIIOI
=
BFMA1lll
&
BFMA1O0l
;
BFMA1lIIOI
=
BFMA1IO0
&
BFMA1O0l
;
BFMA1IlIOI
=
(
BFMA1IIIOI
===
BFMA1lIIOI
)
;
end
if
(
BFMA1l1l
==
1
'b
1
)
begin
BFMA1IIIOI
=
BFMA1OIl
&
BFMA1IIl
;
BFMA1lIIOI
=
GP_IN
&
BFMA1IIl
;
BFMA1llIOI
=
(
BFMA1IIIOI
===
BFMA1lIIOI
)
;
end
BFMA1IOlOI
=
BFMA1I001
|
BFMA1I101
|
BFMA1l001
|
BFMA1O101
|
BFMA1l101
|
BFMA1IO11
|
BFMA1lO11
|
to_boolean
(
BFMA1IlI
|
BFMA1OlI
|
BFMA1lII
|
BFMA1III
|
BFMA1O1l
|
BFMA1I1l
|
BFMA1l1l
)
;
if
(
BFMA1O001
)
begin
case
(
BFMA1IO01
)
BFMA1lI0I
:
begin
if
(
~
BFMA1IOlOI
)
begin
if
(
BFMA1lI11
<=
1
)
begin
BFMA1O001
=
0
;
end
else
begin
BFMA1lI11
=
BFMA1lI11
-
1
;
end
end
end
BFMA1OO0I
:
begin
if
(
BFMA1lI11
<=
1
)
begin
BFMA1O001
=
0
;
end
else
begin
BFMA1lI11
=
BFMA1lI11
-
1
;
end
end
BFMA1l1Ol
,
BFMA1OOIl
:
begin
if
(
$time
>=
BFMA1O00OI
)
begin
BFMA1O001
=
0
;
end
end
BFMA1I1II
,
BFMA1O1II
,
BFMA1l0II
:
begin
if
(
BFMA1IlOOI
==
256
)
begin
BFMA1I1lOI
=
(
INTERRUPT
!=
BFMA1Ol1
)
;
end
else
begin
BFMA1I1lOI
=
(
(
INTERRUPT
[
BFMA1IlOOI
]
)
===
1
'b
1
)
;
end
if
(
BFMA1I1lOI
)
begin
if
(
DEBUG
>=
2
)
$display
(
"BFM:Interrupt Wait Time %0d cycles"
,
BFMA1OOIOI
)
;
BFMA1O001
=
0
;
end
end
BFMA1OOlI
:
begin
BFMA1OI0
<=
BFMA1Ol01
;
BFMA1lO0
<=
BFMA1Il01
;
BFMA1l0l
<=
1
'b
1
;
BFMA1O001
=
0
;
end
BFMA1lIlI
:
begin
BFMA1OI0
<=
BFMA1l011
+
BFMA1I111
;
BFMA1lO0
<=
BFMA1OOOOI
[
BFMA1I111
]
;
BFMA1l0l
<=
1
'b
1
;
BFMA1I111
=
BFMA1I111
+
1
;
if
(
BFMA1I111
>=
BFMA1O111
)
begin
BFMA1O001
=
0
;
end
end
BFMA1IOlI
,
BFMA1lOlI
,
BFMA1OIlI
:
begin
BFMA1OI0
<=
BFMA1Ol01
;
BFMA1OIl
<=
BFMA1Il01
;
BFMA1IIl
<=
BFMA1ll01
;
BFMA1lIl
<=
BFMA1l01
;
BFMA1Oll
<=
1
'b
1
;
if
(
BFMA1I1l
==
1
'b
1
)
begin
BFMA1O001
=
0
;
end
end
BFMA1IIlI
:
begin
if
(
EXT_WAIT
==
1
'b
0
&
BFMA1lI11
==
0
)
begin
if
(
DEBUG
>=
2
)
$display
(
"BFM:Exteral Wait Time %0d cycles"
,
BFMA1OOIOI
)
;
BFMA1O001
=
0
;
end
if
(
BFMA1lI11
>=
1
)
begin
BFMA1lI11
=
BFMA1lI11
-
1
;
end
end
BFMA1IlII
,
BFMA1llII
,
BFMA1l1OI
,
BFMA1OlII
:
begin
BFMA1Oll
<=
1
'b
1
;
BFMA1OIl
<=
BFMA1Il01
;
BFMA1IIl
<=
BFMA1ll01
;
BFMA1lIl
<=
BFMA1l01
;
BFMA1O001
=
0
;
end
BFMA1OOII
:
begin
BFMA1OIl
<=
BFMA1Il01
;
BFMA1IIl
<=
BFMA1ll01
;
BFMA1lIl
<=
BFMA1l01
;
BFMA1l1l
<=
1
'b
1
;
BFMA1Oll
<=
1
'b
0
;
if
(
BFMA1l1l
==
1
'b
1
&
BFMA1llIOI
)
begin
BFMA1l1l
<=
1
'b
0
;
BFMA1O001
=
0
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:GP IO Wait Time %0d cycles"
,
BFMA1OOIOI
)
;
end
end
BFMA1O00I
,
BFMA1I00I
:
begin
case
(
BFMA1lOO1
)
BFMA1Ol10
:
BFMA1O001
=
0
;
BFMA1Il10
:
begin
BFMA1OlO1
=
BFMA1lI
[
1
]
+
BFMA1lI
[
2
]
;
BFMA1I110
=
BFMA1lI
[
3
]
;
BFMA1l110
=
BFMA1lI
[
4
]
%
65536
;
BFMA1IOI1
=
(
(
BFMA1lll1
[
4
]
[
16
]
)
==
1
'b
1
)
;
BFMA1lOI1
=
(
(
BFMA1lll1
[
4
]
[
17
]
)
==
1
'b
1
)
;
BFMA1OII1
=
(
(
BFMA1lll1
[
4
]
[
18
]
)
==
1
'b
1
)
;
BFMA1OOO1
=
BFMA1lI
[
5
]
;
BFMA1IOO1
=
BFMA1lI
[
6
]
;
if
(
~
BFMA1OII1
)
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<
MAX_MEMTEST
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
BFMA1OIO1
[
BFMA1I0I0
]
=
0
;
BFMA1O0O1
=
0
;
BFMA1I0O1
=
0
;
BFMA1l0O1
=
0
;
BFMA1OOI1
=
0
;
BFMA1III1
=
0
;
if
(
BFMA1IO01
==
BFMA1I00I
)
begin
BFMA1OlO1
=
BFMA1lI
[
1
]
;
BFMA1IlO1
=
BFMA1lI
[
2
]
-
BFMA1I110
;
BFMA1I110
=
2
*
BFMA1I110
;
BFMA1OOI1
=
1
;
end
if
(
BFMA1IO01
==
BFMA1O00I
)
begin
$display
(
"BFM:%0d: memtest Started at %0d ns"
,
BFMA1l01
,
$time
)
;
$display
(
"BFM:  Address %08x Size %0d Cycles %5d"
,
BFMA1OlO1
,
BFMA1I110
,
BFMA1OOO1
)
;
end
else
begin
$display
(
"BFM:%0d: dual memtest Started at %0d ns"
,
BFMA1l01
,
$time
)
;
$display
(
"BFM:  Address %08x %08x  Size %0d Cycles %5d"
,
BFMA1OlO1
,
BFMA1IlO1
+
BFMA1I110
/
2
,
BFMA1I110
/
2
,
BFMA1OOO1
)
;
end
case
(
BFMA1l110
)
0
:
begin
end
1
:
$display
(
"BFM: Transfers are APB Byte aligned"
)
;
2
:
$display
(
"BFM: Transfers are APB Half Word aligned"
)
;
3
:
$display
(
"BFM: Transfers are APB Word aligned"
)
;
4
:
$display
(
"BFM: Byte Writes Suppressed"
)
;
default
:
$display
(
"Illegal Align on memtest (FAILURE)"
)
;
endcase
if
(
BFMA1OII1
)
begin
$display
(
"BFM: memtest restarted"
)
;
end
if
(
BFMA1IOI1
)
begin
$display
(
"BFM: Memtest Filling Memory"
)
;
BFMA1lOO1
=
BFMA1I010
;
end
else
if
(
BFMA1OOO1
>
0
)
begin
$display
(
"BFM: Memtest Random Read Writes"
)
;
BFMA1lOO1
=
BFMA1ll10
;
end
else
if
(
BFMA1lOI1
)
begin
$display
(
"BFM: Memtest Verifying Memory Content"
)
;
BFMA1lOO1
=
BFMA1l010
;
end
else
begin
BFMA1lOO1
=
BFMA1O010
;
end
end
BFMA1ll10
,
BFMA1I010
,
BFMA1l010
:
begin
if
(
~
(
BFMA1I101
|
BFMA1I001
)
)
begin
case
(
BFMA1lOO1
)
BFMA1ll10
:
begin
BFMA1IOO1
=
BFMA1lIl0
(
BFMA1IOO1
)
;
BFMA1IIO1
=
BFMA1O1l0
(
BFMA1IOO1
,
BFMA1I110
)
;
BFMA1IOO1
=
BFMA1lIl0
(
BFMA1IOO1
)
;
BFMA1lIO1
=
BFMA1O1l0
(
BFMA1IOO1
,
8
)
;
end
BFMA1I010
:
begin
BFMA1IIO1
=
BFMA1III1
;
BFMA1lIO1
=
6
;
end
BFMA1l010
:
begin
BFMA1IIO1
=
BFMA1III1
;
BFMA1lIO1
=
2
;
end
default
:
begin
end
endcase
case
(
BFMA1l110
)
0
:
begin
end
1
:
begin
BFMA1IIO1
=
4
*
(
BFMA1IIO1
/
4
)
;
case
(
BFMA1lIO1
)
0
,
4
:
begin
BFMA1lIO1
=
BFMA1lIO1
;
end
1
,
5
:
begin
BFMA1lIO1
=
BFMA1lIO1
-
1
;
end
2
,
6
:
begin
BFMA1lIO1
=
BFMA1lIO1
-
2
;
end
default
:
begin
end
endcase
end
2
:
begin
BFMA1IIO1
=
4
*
(
BFMA1IIO1
/
4
)
;
case
(
BFMA1lIO1
)
0
,
4
:
begin
BFMA1lIO1
=
BFMA1lIO1
+
1
;
end
1
,
5
:
begin
BFMA1lIO1
=
BFMA1lIO1
;
end
2
,
6
:
begin
BFMA1lIO1
=
BFMA1lIO1
-
1
;
end
default
:
begin
end
endcase
end
3
:
begin
BFMA1IIO1
=
4
*
(
BFMA1IIO1
/
4
)
;
case
(
BFMA1lIO1
)
0
,
4
:
begin
BFMA1lIO1
=
BFMA1lIO1
+
2
;
end
1
,
5
:
begin
BFMA1lIO1
=
BFMA1lIO1
+
1
;
end
2
,
6
:
begin
BFMA1lIO1
=
BFMA1lIO1
;
end
default
:
begin
end
endcase
end
4
:
begin
case
(
BFMA1lIO1
)
4
:
begin
BFMA1IIO1
=
2
*
(
BFMA1IIO1
/
2
)
;
BFMA1lIO1
=
5
;
end
default
:
begin
end
endcase
end
default
:
begin
end
endcase
if
(
BFMA1lIO1
>=
0
&
BFMA1lIO1
<=
2
)
begin
case
(
BFMA1lIO1
)
0
:
begin
BFMA1lI01
=
3
'b
000
;
BFMA1IIO1
=
BFMA1IIO1
;
BFMA1llO1
=
(
BFMA1OIO1
[
BFMA1IIO1
+
0
]
>=
256
)
;
end
1
:
begin
BFMA1lI01
=
3
'b
001
;
BFMA1IIO1
=
2
*
(
BFMA1IIO1
/
2
)
;
BFMA1llO1
=
(
(
BFMA1OIO1
[
BFMA1IIO1
+
0
]
>=
256
)
&
(
BFMA1OIO1
[
BFMA1IIO1
+
1
]
>=
256
)
)
;
end
2
:
begin
BFMA1lI01
=
3
'b
010
;
BFMA1IIO1
=
4
*
(
BFMA1IIO1
/
4
)
;
BFMA1llO1
=
(
(
BFMA1OIO1
[
BFMA1IIO1
+
0
]
>=
256
)
&
(
BFMA1OIO1
[
BFMA1IIO1
+
1
]
>=
256
)
&
(
BFMA1OIO1
[
BFMA1IIO1
+
2
]
>=
256
)
&
(
BFMA1OIO1
[
BFMA1IIO1
+
3
]
>=
256
)
)
;
end
default
:
begin
end
endcase
if
(
BFMA1llO1
)
begin
BFMA1I001
=
1
;
BFMA1O0O1
=
BFMA1O0O1
+
1
;
if
(
BFMA1OOI1
==
1
&
BFMA1IIO1
>=
BFMA1I110
/
2
)
begin
BFMA1Ol01
=
BFMA1IlO1
+
BFMA1IIO1
;
end
else
begin
BFMA1Ol01
=
BFMA1OlO1
+
BFMA1IIO1
;
end
case
(
BFMA1lIO1
)
0
:
begin
BFMA1Il01
=
{
BFMA1lI1
[
31
:
8
]
,
BFMA1OIO1
[
BFMA1IIO1
+
0
]
[
7
:
0
]
}
;
end
1
:
begin
BFMA1Il01
=
{
BFMA1lI1
[
31
:
16
]
,
BFMA1OIO1
[
BFMA1IIO1
+
1
]
[
7
:
0
]
,
BFMA1OIO1
[
BFMA1IIO1
+
0
]
[
7
:
0
]
}
;
end
2
:
begin
BFMA1Il01
=
{
BFMA1OIO1
[
BFMA1IIO1
+
3
]
[
7
:
0
]
,
BFMA1OIO1
[
BFMA1IIO1
+
2
]
[
7
:
0
]
,
BFMA1OIO1
[
BFMA1IIO1
+
1
]
[
7
:
0
]
,
BFMA1OIO1
[
BFMA1IIO1
+
0
]
[
7
:
0
]
}
;
end
default
:
begin
BFMA1Il01
=
BFMA1lI1
[
31
:
0
]
;
end
endcase
BFMA1ll01
=
{
32
{
1
'b
1
}
}
;
end
else
begin
BFMA1lIO1
=
BFMA1lIO1
+
4
;
if
(
BFMA1lIO1
==
4
&
BFMA1l110
==
4
)
begin
BFMA1lIO1
=
5
;
end
end
end
if
(
BFMA1lIO1
>=
4
&
BFMA1lIO1
<=
6
)
begin
BFMA1I101
=
1
;
BFMA1I0O1
=
BFMA1I0O1
+
1
;
BFMA1IOO1
=
BFMA1lIl0
(
BFMA1IOO1
)
;
BFMA1Il01
=
BFMA1IOO1
;
case
(
BFMA1lIO1
)
4
:
begin
BFMA1lI01
=
3
'b
000
;
BFMA1IIO1
=
BFMA1IIO1
;
BFMA1OIO1
[
BFMA1IIO1
+
0
]
=
256
+
BFMA1Il01
[
7
:
0
]
;
end
5
:
begin
BFMA1lI01
=
3
'b
001
;
BFMA1IIO1
=
2
*
(
BFMA1IIO1
/
2
)
;
BFMA1OIO1
[
BFMA1IIO1
+
0
]
=
256
+
BFMA1Il01
[
7
:
0
]
;
BFMA1OIO1
[
BFMA1IIO1
+
1
]
=
256
+
BFMA1Il01
[
15
:
8
]
;
end
6
:
begin
BFMA1lI01
=
3
'b
010
;
BFMA1IIO1
=
4
*
(
BFMA1IIO1
/
4
)
;
BFMA1OIO1
[
BFMA1IIO1
+
0
]
=
256
+
BFMA1Il01
[
7
:
0
]
;
BFMA1OIO1
[
BFMA1IIO1
+
1
]
=
256
+
BFMA1Il01
[
15
:
8
]
;
BFMA1OIO1
[
BFMA1IIO1
+
2
]
=
256
+
BFMA1Il01
[
23
:
16
]
;
BFMA1OIO1
[
BFMA1IIO1
+
3
]
=
256
+
BFMA1Il01
[
31
:
24
]
;
end
default
:
begin
end
endcase
if
(
BFMA1OOI1
==
1
&
BFMA1IIO1
>=
BFMA1I110
/
2
)
begin
BFMA1Ol01
=
BFMA1IlO1
+
BFMA1IIO1
;
end
else
begin
BFMA1Ol01
=
BFMA1OlO1
+
BFMA1IIO1
;
end
end
if
(
BFMA1lIO1
==
3
|
BFMA1lIO1
==
7
)
begin
BFMA1l0O1
=
BFMA1l0O1
+
1
;
end
BFMA1III1
=
BFMA1III1
+
4
;
case
(
BFMA1lOO1
)
BFMA1ll10
:
begin
if
(
BFMA1OOO1
>
0
)
begin
BFMA1OOO1
=
BFMA1OOO1
-
1
;
end
else
if
(
BFMA1lOI1
)
begin
BFMA1III1
=
0
;
BFMA1lOO1
=
BFMA1l010
;
$display
(
"BFM: Memtest Verifying Memory Content"
)
;
end
else
begin
BFMA1lOO1
=
BFMA1O010
;
end
end
BFMA1I010
:
begin
if
(
BFMA1III1
>=
BFMA1I110
)
begin
if
(
BFMA1OOO1
==
0
)
begin
if
(
BFMA1lOI1
)
begin
BFMA1III1
=
0
;
BFMA1lOO1
=
BFMA1l010
;
$display
(
"BFM: Memtest Verifying Memory Content"
)
;
end
else
begin
BFMA1lOO1
=
BFMA1O010
;
end
end
else
begin
BFMA1lOO1
=
BFMA1ll10
;
$display
(
"BFM: Memtest Random Read Writes"
)
;
end
end
end
BFMA1l010
:
begin
if
(
BFMA1III1
>=
BFMA1I110
)
begin
BFMA1lOO1
=
BFMA1O010
;
end
end
default
:
begin
end
endcase
BFMA1Il11
=
BFMA1II01
;
end
end
BFMA1O010
:
begin
if
(
~
BFMA1IOlOI
)
begin
BFMA1lOO1
=
BFMA1Ol10
;
$display
(
"BFM: bfmtest complete  Writes %0d  Reads %0d  Nops %0d"
,
BFMA1I0O1
,
BFMA1O0O1
,
BFMA1l0O1
)
;
end
end
endcase
end
default
:
begin
end
endcase
end
if
(
BFMA1OO0OI
==
0
)
begin
BFMA1IO0OI
=
0
;
BFMA1OO0OI
=
BFMA1IllOI
;
end
else
begin
BFMA1OO0OI
=
BFMA1OO0OI
-
1
;
BFMA1IO0OI
=
1
;
end
if
(
HREADY
==
1
'b
1
)
begin
BFMA1l0
<=
2
'b
00
;
BFMA1O1
<=
1
'b
0
;
BFMA1lII
<=
1
'b
0
;
BFMA1OlI
<=
1
'b
0
;
BFMA1llI
<=
1
'b
0
;
if
(
BFMA1lII
==
1
'b
1
|
BFMA1OlI
==
1
'b
1
)
begin
BFMA1I0I
<=
1
'b
0
;
end
if
(
BFMA1I101
&
HREADY
==
1
'b
1
)
begin
BFMA1l1
<=
BFMA1Ol01
;
BFMA1O1
<=
1
'b
1
;
BFMA1ll
<=
BFMA1l1IOI
;
BFMA1l0
<=
2
'b
10
;
BFMA1O0
<=
BFMA1O1IOI
;
BFMA1I0
<=
BFMA1I1IOI
;
BFMA1IOI
<=
BFMA1lI01
;
BFMA1l1I
<=
BFMA1l01l
(
BFMA1lI01
,
BFMA1Ol01
[
1
:
0
]
,
BFMA1Il01
,
BFMA1I0lOI
)
;
BFMA1lII
<=
1
'b
1
;
BFMA1O00
<=
BFMA1l01
;
BFMA1I101
=
0
;
end
if
(
BFMA1I001
&
HREADY
==
1
'b
1
)
begin
BFMA1l1
<=
BFMA1Ol01
;
BFMA1O1
<=
1
'b
0
;
BFMA1ll
<=
BFMA1l1IOI
;
BFMA1l0
<=
2
'b
10
;
BFMA1O0
<=
BFMA1O1IOI
;
BFMA1I0
<=
BFMA1I1IOI
;
BFMA1IOI
<=
BFMA1lI01
;
BFMA1O1I
<=
BFMA1l01l
(
BFMA1lI01
,
BFMA1Ol01
[
1
:
0
]
,
BFMA1Il01
,
BFMA1I0lOI
)
;
BFMA1I1I
<=
BFMA1OIO0
(
BFMA1lI01
,
BFMA1Ol01
[
1
:
0
]
,
BFMA1ll01
,
BFMA1I0lOI
)
;
BFMA1O00
<=
BFMA1l01
;
BFMA1OlI
<=
1
'b
1
;
BFMA1I0I
<=
1
'b
1
;
BFMA1I001
=
0
;
end
if
(
BFMA1IO11
&
HREADY
==
1
'b
1
)
begin
BFMA1l1
<=
BFMA1Ol01
;
BFMA1O1
<=
BFMA1I00OI
;
BFMA1ll
<=
BFMA1I10OI
;
BFMA1l0
<=
BFMA1l00OI
;
BFMA1O0
<=
BFMA1l10OI
;
BFMA1I0
<=
BFMA1O10OI
;
BFMA1IOI
<=
BFMA1lI01
;
BFMA1l1I
<=
BFMA1l01l
(
BFMA1lI01
,
BFMA1Ol01
[
1
:
0
]
,
BFMA1Il01
,
BFMA1I0lOI
)
;
BFMA1lII
<=
1
'b
1
;
BFMA1O00
<=
BFMA1l01
;
BFMA1IO11
=
0
;
end
if
(
BFMA1l101
&
HREADY
==
1
'b
1
)
begin
BFMA1l1
<=
BFMA1Ol01
;
BFMA1O1
<=
1
'b
0
;
BFMA1ll
<=
BFMA1l1IOI
;
BFMA1O0
<=
BFMA1O1IOI
;
BFMA1I0
<=
BFMA1I1IOI
;
BFMA1IOI
<=
BFMA1lI01
;
BFMA1O1I
<=
BFMA1l01l
(
BFMA1lI01
,
BFMA1Ol01
[
1
:
0
]
,
BFMA1Il01
,
BFMA1I0lOI
)
;
BFMA1I1I
<=
BFMA1OIO0
(
BFMA1lI01
,
BFMA1Ol01
[
1
:
0
]
,
BFMA1ll01
,
BFMA1I0lOI
)
;
BFMA1O00
<=
BFMA1l01
;
if
(
BFMA1OlI
==
1
'b
1
|
BFMA1IlI
==
1
'b
1
)
begin
BFMA1l0
<=
2
'b
00
;
end
else
begin
BFMA1l0
<=
2
'b
10
;
BFMA1OlI
<=
1
'b
1
;
BFMA1llI
<=
1
'b
1
;
end
if
(
BFMA1O0I
==
1
'b
1
&
BFMA1OlIOI
)
begin
BFMA1l101
=
0
;
end
end
if
(
BFMA1l001
&
HREADY
==
1
'b
1
)
begin
BFMA1l1
<=
BFMA1Ol01
;
BFMA1O1
<=
1
'b
1
;
BFMA1ll
<=
BFMA1l1IOI
;
BFMA1O0
<=
BFMA1O1IOI
;
BFMA1I0
<=
BFMA1I1IOI
;
BFMA1IOI
<=
BFMA1lI01
;
BFMA1O00
<=
BFMA1l01
;
if
(
BFMA1IO0OI
)
begin
BFMA1l0
<=
2
'b
01
;
end
else
begin
BFMA1l1I
<=
BFMA1l01l
(
BFMA1lI01
,
BFMA1Ol01
[
1
:
0
]
,
to_slv32
(
BFMA1OOOOI
[
BFMA1I111
]
)
,
BFMA1I0lOI
)
;
BFMA1lII
<=
1
'b
1
;
if
(
BFMA1I111
==
0
|
BFMA1l1l1
==
3
|
bound1k
(
BFMA1O0lOI
,
BFMA1Ol01
)
)
begin
BFMA1l0
<=
2
'b
10
;
end
else
begin
BFMA1l0
<=
2
'b
11
;
end
BFMA1Ol01
=
BFMA1Ol01
+
BFMA1l111
;
BFMA1I111
=
BFMA1I111
+
1
;
if
(
BFMA1I111
==
BFMA1O111
)
begin
BFMA1l001
=
0
;
end
end
end
if
(
BFMA1O101
&
HREADY
==
1
'b
1
)
begin
BFMA1l1
<=
BFMA1Ol01
;
BFMA1O1
<=
1
'b
0
;
BFMA1ll
<=
BFMA1l1IOI
;
BFMA1O0
<=
BFMA1O1IOI
;
BFMA1I0
<=
BFMA1I1IOI
;
BFMA1IOI
<=
BFMA1lI01
;
BFMA1O00
<=
BFMA1l01
;
if
(
BFMA1IO0OI
)
begin
BFMA1l0
<=
2
'b
01
;
end
else
begin
BFMA1O1I
<=
BFMA1l01l
(
BFMA1lI01
,
BFMA1Ol01
[
1
:
0
]
,
to_slv32
(
BFMA1OOOOI
[
BFMA1I111
]
)
,
BFMA1I0lOI
)
;
BFMA1I1I
<=
BFMA1OIO0
(
BFMA1lI01
,
BFMA1Ol01
[
1
:
0
]
,
BFMA1ll01
,
BFMA1I0lOI
)
;
BFMA1OlI
<=
1
'b
1
;
BFMA1I0I
<=
1
'b
1
;
if
(
BFMA1I111
==
0
|
BFMA1l1l1
==
3
|
bound1k
(
BFMA1O0lOI
,
BFMA1Ol01
)
)
begin
BFMA1l0
<=
2
'b
10
;
end
else
begin
BFMA1l0
<=
2
'b
11
;
end
BFMA1Ol01
=
BFMA1Ol01
+
BFMA1l111
;
BFMA1I111
=
BFMA1I111
+
1
;
if
(
BFMA1I111
==
BFMA1O111
)
begin
BFMA1O101
=
0
;
end
end
end
end
if
(
HREADY
==
1
'b
1
)
begin
BFMA1III
<=
BFMA1lII
;
BFMA1IlI
<=
BFMA1OlI
;
BFMA1O0I
<=
BFMA1llI
;
BFMA1l0I
<=
BFMA1I0I
;
BFMA1OOl
<=
BFMA1O1I
;
BFMA1IOl
<=
BFMA1I1I
;
BFMA1I00
<=
BFMA1O00
;
BFMA1OOI
<=
BFMA1l1
;
BFMA1lOI
<=
BFMA1IOI
;
end
BFMA1I1l
<=
BFMA1O1l
;
BFMA1II0
<=
BFMA1OI0
;
BFMA1Ill
<=
BFMA1Oll
;
BFMA1lll
<=
BFMA1OIl
;
BFMA1O0l
<=
BFMA1IIl
;
BFMA1I0l
<=
BFMA1lIl
;
if
(
HREADY
==
1
'b
1
)
begin
if
(
BFMA1lII
==
1
'b
1
)
begin
BFMA1lOl
<=
BFMA1l1I
;
end
else
begin
BFMA1lOl
<=
{
32
{
1
'b
0
}
}
;
end
if
(
BFMA1III
==
1
'b
1
&
DEBUG
>=
3
)
begin
$display
(
"BFM: Data Write %08x %08x"
,
BFMA1OOI
,
BFMA1lOl
)
;
end
if
(
BFMA1lO0OI
&
BFMA1III
==
1
'b
1
)
begin
$fdisplay
(
BFMA1lIl1
,
"%05d AW %c %08x %08x"
,
$time
,
BFMA1IlO0
(
BFMA1lOI
)
,
BFMA1OOI
,
BFMA1lOl
)
;
end
end
if
(
BFMA1OO0
==
1
'b
1
&
BFMA1II0OI
)
begin
$fdisplay
(
BFMA1lIl1
,
"%05d GW   %08x "
,
$time
,
BFMA1O10
)
;
end
if
(
BFMA1l0l
==
1
'b
1
&
BFMA1OI0OI
)
begin
$fdisplay
(
BFMA1lIl1
,
"%05d EW   %08x %08x"
,
$time
,
BFMA1OI0
,
BFMA1lO0
)
;
end
if
(
HREADY
==
1
'b
1
)
begin
if
(
BFMA1IlI
==
1
'b
1
)
begin
if
(
DEBUG
>=
3
)
begin
if
(
BFMA1IOl
==
BFMA1lI1
)
begin
$display
(
"BFM: Data Read %08x %08x"
,
BFMA1OOI
,
HRDATA
)
;
end
else
begin
$display
(
"BFM: Data Read %08x %08x MASK:%08x"
,
BFMA1OOI
,
HRDATA
,
BFMA1IOl
)
;
end
end
if
(
BFMA1lO0OI
)
begin
$fdisplay
(
BFMA1lIl1
,
"%05d AR %c %08x %08x"
,
$time
,
BFMA1IlO0
(
BFMA1lOI
)
,
BFMA1OOI
,
HRDATA
)
;
end
if
(
BFMA1OOlOI
>=
0
)
begin
BFMA1ll1
[
BFMA1OOlOI
]
=
BFMA1O01l
(
BFMA1IIO0
(
BFMA1lOI
,
BFMA1OOI
[
1
:
0
]
,
HRDATA
,
BFMA1I0lOI
)
)
;
end
if
(
BFMA1l0I
==
1
'b
1
&
~
BFMA1OlIOI
)
begin
BFMA1II10
=
BFMA1II10
+
1
;
$display
(
"ERROR: AHB Data Read Comparison failed Addr:%08x  Got:%08x  EXP:%08x  (MASK:%08x)"
,
BFMA1OOI
,
HRDATA
,
BFMA1OOl
,
BFMA1IOl
)
;
$display
(
"       Stimulus file %0s  Line No %0d"
,
BFMA1lOlOI
[
BFMA1OIl0
(
BFMA1I00
,
BFMA1IIlOI
)
]
,
BFMA1l1I0
(
BFMA1I00
,
BFMA1IIlOI
)
)
;
$display
(
"BFM Data Compare Error (ERROR)"
)
;
$stop
;
if
(
BFMA1lO0OI
)
begin
$fdisplay
(
BFMA1lIl1
,
"%05d ERROR  Addr:%08x  Got:%08x  EXP:%08x  (MASK:%08x)"
,
$time
,
BFMA1OOI
,
HRDATA
,
BFMA1OOl
,
BFMA1IOl
)
;
end
end
end
end
if
(
BFMA1l1l
==
1
'b
1
)
begin
if
(
DEBUG
>=
3
)
begin
if
(
BFMA1IIl
==
BFMA1lI1
)
begin
$display
(
"BFM: GP IO Data Read %08x"
,
GP_IN
)
;
end
else
begin
$display
(
"BFM: GP IO Data Read %08x  MASK:%08x"
,
GP_IN
,
BFMA1IIl
)
;
end
end
if
(
BFMA1II0OI
)
begin
$fdisplay
(
BFMA1lIl1
,
"%05d GR   %08x "
,
$time
,
BFMA1OIl
)
;
end
if
(
BFMA1OOlOI
>=
0
)
begin
BFMA1ll1
[
BFMA1OOlOI
]
=
GP_IN
;
end
if
(
BFMA1Oll
==
1
'b
1
&
~
BFMA1llIOI
)
begin
BFMA1II10
=
BFMA1II10
+
1
;
$display
(
"GPIO input not as expected  Got:%08x  EXP:%08x  (MASK:%08x)"
,
GP_IN
,
BFMA1OIl
,
BFMA1IIl
)
;
$display
(
"       Stimulus file %0s  Line No %0d"
,
BFMA1lOlOI
[
BFMA1OIl0
(
BFMA1lIl
,
BFMA1IIlOI
)
]
,
BFMA1l1I0
(
BFMA1lIl
,
BFMA1IIlOI
)
)
;
$display
(
"BFM GPIO Compare Error (ERROR)"
)
;
$stop
;
if
(
BFMA1II0OI
)
begin
$fdisplay
(
BFMA1lIl1
,
"ERROR  Got:%08x  EXP:%08x  (MASK:%08x)"
,
GP_IN
,
BFMA1OIl
,
BFMA1IIl
)
;
end
end
end
if
(
BFMA1I1l
==
1
'b
1
)
begin
if
(
DEBUG
>=
3
)
begin
if
(
BFMA1O0l
==
BFMA1lI1
)
begin
$display
(
"BFM: Extention Data Read %08x %08x"
,
BFMA1II0
,
BFMA1IO0
)
;
end
else
begin
$display
(
"BFM: Extention Data Read %08x %08x  MASK:%08x"
,
BFMA1II0
,
BFMA1IO0
,
BFMA1O0l
)
;
end
end
if
(
BFMA1OI0OI
)
begin
$fdisplay
(
BFMA1lIl1
,
"%05d ER   %08x %08x"
,
$time
,
BFMA1II0
,
BFMA1lll
)
;
end
if
(
BFMA1OOlOI
>=
0
)
begin
BFMA1ll1
[
BFMA1OOlOI
]
=
BFMA1O01l
(
BFMA1IO0
)
;
end
if
(
BFMA1Ill
==
1
'b
1
&
~
BFMA1IlIOI
)
begin
BFMA1II10
=
BFMA1II10
+
1
;
$display
(
"ERROR: Extention Data Read Comparison FAILED  Got:%08x  EXP:%08x  (MASK:%08x)"
,
BFMA1IO0
,
BFMA1lll
,
BFMA1O0l
)
;
$display
(
"       Stimulus file %0s  Line No %0d"
,
BFMA1lOlOI
[
BFMA1OIl0
(
BFMA1I0l
,
BFMA1IIlOI
)
]
,
BFMA1l1I0
(
BFMA1I0l
,
BFMA1IIlOI
)
)
;
$display
(
"BFM Extention Data Compare Error (ERROR)"
)
;
$stop
;
if
(
BFMA1OI0OI
)
begin
$fdisplay
(
BFMA1lIl1
,
"ERROR  Got:%08x  EXP:%08x  (MASK:%08x)"
,
BFMA1IO0
,
BFMA1lll
,
BFMA1O0l
)
;
end
end
end
BFMA1OO1OI
=
BFMA1I001
|
BFMA1I101
|
BFMA1l001
|
BFMA1O101
|
BFMA1l101
|
BFMA1IO11
|
to_boolean
(
BFMA1OlI
|
BFMA1lII
|
BFMA1O1l
|
BFMA1l1l
)
|
(
to_boolean
(
(
BFMA1IlI
|
BFMA1III
)
&
~
HREADY
)
)
;
if
(
BFMA1O001
)
begin
case
(
BFMA1IO01
)
BFMA1OI1I
:
begin
if
(
~
BFMA1OO1OI
)
begin
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:checktime was %0d cycles "
,
BFMA1l01
,
BFMA1OOIOI
)
;
if
(
BFMA1OOIOI
<
BFMA1lI
[
1
]
|
BFMA1OOIOI
>
BFMA1lI
[
2
]
)
begin
$display
(
"BFM: ERROR checktime %0d %0d Actual %0d"
,
BFMA1lI
[
1
]
,
BFMA1lI
[
2
]
,
BFMA1OOIOI
)
;
$display
(
"       Stimulus file %0s  Line No %0d"
,
BFMA1lOlOI
[
BFMA1OIl0
(
BFMA1I00
,
BFMA1IIlOI
)
]
,
BFMA1l1I0
(
BFMA1I00
,
BFMA1IIlOI
)
)
;
$display
(
"BFM checktime failure (ERROR)"
)
;
BFMA1II10
=
BFMA1II10
+
1
;
$stop
;
end
BFMA1O001
=
0
;
BFMA1I1O1
=
BFMA1OOIOI
;
end
end
BFMA1Ol1I
:
begin
if
(
~
BFMA1OO1OI
)
begin
BFMA1l1O1
=
BFMA1l1O1
-
1
;
if
(
DEBUG
>=
2
)
$display
(
"BFM:%0d:checktimer was %0d cycles "
,
BFMA1l01
,
BFMA1l1O1
)
;
if
(
BFMA1l1O1
<
BFMA1lI
[
1
]
|
BFMA1l1O1
>
BFMA1lI
[
2
]
)
begin
$display
(
"BFM: ERROR checktimer %0d %0d Actual %0d"
,
BFMA1lI
[
1
]
,
BFMA1lI
[
2
]
,
BFMA1l1O1
)
;
$display
(
"       Stimulus file %0s  Line No %0d"
,
BFMA1lOlOI
[
BFMA1OIl0
(
BFMA1I00
,
BFMA1IIlOI
)
]
,
BFMA1l1I0
(
BFMA1I00
,
BFMA1IIlOI
)
)
;
$display
(
"BFM checktimer failure (ERROR)"
)
;
BFMA1II10
=
BFMA1II10
+
1
;
$stop
;
end
BFMA1O001
=
0
;
BFMA1O1O1
=
BFMA1l1O1
;
end
end
default
:
begin
end
endcase
end
if
(
BFMA1l0lOI
)
begin
if
(
BFMA1Il11
>
0
)
begin
BFMA1Il11
=
BFMA1Il11
-
1
;
end
else
begin
BFMA1Il11
=
BFMA1II01
;
$display
(
"BFM Command Timeout Occured"
)
;
$display
(
"       Stimulus file %0s  Line No %0d"
,
BFMA1lOlOI
[
BFMA1OIl0
(
BFMA1I00
,
BFMA1IIlOI
)
]
,
BFMA1l1I0
(
BFMA1I00
,
BFMA1IIlOI
)
)
;
if
(
~
BFMA1lOOOI
)
$display
(
"BFM Command timeout occured (ERROR)"
)
;
if
(
BFMA1lOOOI
)
$display
(
"BFM Completed and timeout occured (ERROR)"
)
;
$stop
;
end
end
else
begin
BFMA1Il11
=
BFMA1II01
;
end
if
(
BFMA1II10
>
0
)
begin
BFMA1OO1
<=
1
'b
1
;
end
if
(
BFMA1O001
|
BFMA1I001
|
BFMA1I101
|
BFMA1l001
|
BFMA1O101
|
BFMA1l101
|
BFMA1IO11
|
(
(
BFMA1OO11
|
BFMA1lllOI
)
&
BFMA1IOlOI
)
)
begin
BFMA1OI11
=
1
;
end
else
begin
BFMA1OO11
=
0
;
if
(
~
BFMA1lOOOI
)
begin
BFMA1OI11
=
0
;
end
BFMA1O000
=
BFMA1O000
+
BFMA1OI01
;
BFMA1OI01
=
0
;
if
(
OPMODE
>
0
)
begin
if
(
BFMA1O1lOI
|
BFMA1lOOOI
)
begin
BFMA1l0lOI
=
0
;
BFMA1OI11
=
0
;
end
end
end
if
(
BFMA1l10
==
1
'b
0
&
OPMODE
==
0
&
BFMA1lOOOI
&
~
BFMA1IOlOI
)
begin
$display
(
"###########################################################"
)
;
$display
(
" "
)
;
if
(
BFMA1II10
==
0
)
begin
$display
(
"BFM Simulation Complete - %0d Instructions - NO ERRORS"
,
BFMA1IOIOI
)
;
end
else
begin
$display
(
"BFM Simulation Complete - %0d Instructions - %0d ERRORS OCCURED"
,
BFMA1IOIOI
,
BFMA1II10
)
;
end
$display
(
" "
)
;
$display
(
"###########################################################"
)
;
$display
(
" "
)
;
BFMA1l10
<=
1
'b
1
;
BFMA1OI11
=
1
;
BFMA1l0lOI
=
0
;
if
(
BFMA1O11
)
begin
$fflush
(
BFMA1lIl1
)
;
$fclose
(
BFMA1lIl1
)
;
end
if
(
BFMA1l1lOI
==
1
)
$stop
;
if
(
BFMA1l1lOI
==
2
)
$finish
;
end
CON_BUSY
<=
(
BFMA1l0lOI
|
BFMA1IOlOI
)
;
INSTR_OUT
<=
to_slv32
(
BFMA1O000
)
;
end
end
assign
#
TPD
GP_OUT
=
BFMA1O10
;
assign
#
TPD
EXT_WR
=
BFMA1l0l
;
assign
#
TPD
EXT_RD
=
BFMA1O1l
;
assign
#
TPD
EXT_ADDR
=
BFMA1OI0
;
assign
#
TPD
EXT_DATA
=
(
BFMA1l0l
==
1
'b
1
)
?
BFMA1lO0
:
{
32
{
1
'b
z
}
}
;
assign
BFMA1IO0
=
EXT_DATA
;
always
@
(
BFMA1l1
)
begin
begin
:
BFMA1l0OII
integer
BFMA1I0I0
;
for
(
BFMA1I0I0
=
0
;
BFMA1I0I0
<=
15
;
BFMA1I0I0
=
BFMA1I0I0
+
1
)
begin
BFMA1OII
[
BFMA1I0I0
]
<=
(
BFMA1l1
[
31
:
28
]
==
BFMA1I0I0
)
;
end
end
end
assign
HCLK
=
(
BFMA1IO1
)
?
1
'b
x
:
(
SYSCLK
|
BFMA1l00
)
;
assign
PCLK
=
(
BFMA1IO1
)
?
1
'b
x
:
(
SYSCLK
|
BFMA1l00
)
;
assign
#
TPD
HRESETN
=
(
BFMA1lO1
)
?
1
'b
x
:
BFMA1Il
;
assign
#
TPD
HADDR
=
(
BFMA1OI1
)
?
{
32
{
1
'b
x
}
}
:
BFMA1l1
;
assign
#
TPD
HWDATA
=
(
BFMA1II1
)
?
{
32
{
1
'b
x
}
}
:
BFMA1lOl
;
assign
#
TPD
HBURST
=
(
BFMA1OI1
)
?
{
3
{
1
'b
x
}
}
:
BFMA1ll
;
assign
#
TPD
HMASTLOCK
=
(
BFMA1OI1
)
?
1
'b
x
:
BFMA1O0
;
assign
#
TPD
HPROT
=
(
BFMA1OI1
)
?
{
4
{
1
'b
x
}
}
:
BFMA1I0
;
assign
#
TPD
HSIZE
=
(
BFMA1OI1
)
?
{
3
{
1
'b
x
}
}
:
BFMA1IOI
;
assign
#
TPD
HTRANS
=
(
BFMA1OI1
)
?
{
2
{
1
'b
x
}
}
:
BFMA1l0
;
assign
#
TPD
HWRITE
=
(
BFMA1OI1
)
?
1
'b
x
:
BFMA1O1
;
assign
#
TPD
HSEL
=
(
BFMA1OI1
)
?
{
16
{
1
'b
x
}
}
:
BFMA1OII
;
assign
#
TPD
CON_DATA
=
(
BFMA1Il0
==
1
'b
1
)
?
BFMA1Ol0
:
{
32
{
1
'b
z
}
}
;
assign
BFMA1lI0
=
CON_DATA
;
assign
#
TPD
FINISHED
=
BFMA1l10
;
assign
#
TPD
FAILED
=
BFMA1OO1
;
endmodule
