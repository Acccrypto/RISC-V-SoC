//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Sun Nov 26 17:03:04 2023
// Version: 2022.2 2022.2.0.10
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// MSS_WRAPPER
module MSS_WRAPPER(
    // Inputs
    CAN_0_RXBUS_F2M,
    CAN_1_RXBUS,
    FIC_0_ACLK,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARREADY,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWREADY,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BRESP,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BVALID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RDATA,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RLAST,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RRESP,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RVALID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WREADY,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARADDR,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARBURST,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARCACHE,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLEN,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLOCK,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARPROT,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARQOS,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARSIZE,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARVALID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWADDR,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWBURST,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWCACHE,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLEN,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLOCK,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWPROT,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWQOS,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWSIZE,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWVALID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BREADY,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RREADY,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WDATA,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WLAST,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WSTRB,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WVALID,
    FIC_1_ACLK,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARREADY,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWREADY,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BRESP,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BVALID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RDATA,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RLAST,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RRESP,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RVALID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WREADY,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARADDR,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARBURST,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARCACHE,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLEN,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLOCK,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARPROT,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARQOS,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARSIZE,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARVALID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWADDR,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWBURST,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWCACHE,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLEN,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLOCK,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWPROT,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWQOS,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWSIZE,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWVALID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BREADY,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RREADY,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WDATA,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WLAST,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WSTRB,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WVALID,
    FIC_2_ACLK,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARADDR,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARBURST,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARCACHE,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLEN,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLOCK,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARPROT,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARQOS,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARSIZE,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARVALID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWADDR,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWBURST,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWCACHE,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLEN,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLOCK,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWPROT,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWQOS,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWSIZE,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWVALID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BREADY,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RREADY,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WDATA,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WLAST,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WSTRB,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WVALID,
    FIC_3_APB_INITIATOR_FIC_3_APB_M_PRDATA,
    FIC_3_APB_INITIATOR_FIC_3_APB_M_PREADY,
    FIC_3_APB_INITIATOR_FIC_3_APB_M_PSLVERR,
    FIC_3_PCLK,
    GPIO_2_F2M_30,
    GPIO_2_F2M_31,
    MMUART_0_RXD_F2M,
    MMUART_1_RXD_F2M,
    MMUART_2_RXD_F2M,
    MMUART_3_RXD_F2M,
    MMUART_4_RXD_F2M,
    MSS_INT_F2M_0,
    MSS_INT_F2M_2,
    MSS_INT_F2M_3,
    MSS_RESET_N_F2M,
    REFCLK,
    REFCLK_N,
    SD_CD_EMMC_STRB,
    SD_WP_EMMC_RSTN,
    SGMII_RX0_N,
    SGMII_RX0_P,
    SGMII_RX1_N,
    SGMII_RX1_P,
    SPI_1_DI,
    USB_CLK,
    USB_DIR,
    USB_NXT,
    // Outputs
    CA,
    CAN_0_TXBUS_M2F,
    CAN_0_TX_EBL_M2F,
    CAN_1_TXBUS,
    CAN_1_TX_EBL_N,
    CK,
    CKE,
    CK_N,
    CS,
    DM,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARADDR,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARBURST,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARCACHE,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARLEN,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARLOCK,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARPROT,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARQOS,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARSIZE,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARVALID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWADDR,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWBURST,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWCACHE,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWLEN,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWLOCK,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWPROT,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWQOS,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWSIZE,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWVALID,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BREADY,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RREADY,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WDATA,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WLAST,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WSTRB,
    FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WVALID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARREADY,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWREADY,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BRESP,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BVALID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RDATA,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RLAST,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RRESP,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RVALID,
    FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WREADY,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARADDR,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARBURST,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARCACHE,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARLEN,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARLOCK,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARPROT,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARQOS,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARSIZE,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARVALID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWADDR,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWBURST,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWCACHE,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWLEN,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWLOCK,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWPROT,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWQOS,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWSIZE,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWVALID,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BREADY,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RREADY,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WDATA,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WLAST,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WSTRB,
    FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WVALID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARREADY,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWREADY,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BRESP,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BVALID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RDATA,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RLAST,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RRESP,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RVALID,
    FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WREADY,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARREADY,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWREADY,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BRESP,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BVALID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RDATA,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RLAST,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RRESP,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RVALID,
    FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WREADY,
    FIC_3_APB_INITIATOR_FIC_3_APB_M_PADDR,
    FIC_3_APB_INITIATOR_FIC_3_APB_M_PENABLE,
    FIC_3_APB_INITIATOR_FIC_3_APB_M_PSEL,
    FIC_3_APB_INITIATOR_FIC_3_APB_M_PWDATA,
    FIC_3_APB_INITIATOR_FIC_3_APB_M_PWRITE,
    GPIO_2_M2F_16,
    GPIO_2_M2F_17,
    GPIO_2_M2F_18,
    GPIO_2_M2F_19,
    GPIO_2_M2F_26,
    GPIO_2_M2F_27,
    GPIO_2_M2F_28,
    MAC_1_MDC,
    MMUART_0_TXD_M2F,
    MMUART_1_TXD_M2F,
    MMUART_2_TXD_M2F,
    MMUART_3_TXD_M2F,
    MMUART_4_TXD_M2F,
    MSS_DLL_LOCKS,
    MSS_RESET_N_M2F,
    ODT,
    RESET_N,
    SD_CLK_EMMC_CLK,
    SD_POW_EMMC_DATA4,
    SD_VOLT_CMD_DIR_EMMC_DATA7,
    SD_VOLT_DIR_0_EMMC_UNUSED,
    SD_VOLT_DIR_1_3_EMMC_UNUSED,
    SD_VOLT_EN_EMMC_DATA6,
    SD_VOLT_SEL_EMMC_DATA5,
    SGMII_TX0_N,
    SGMII_TX0_P,
    SGMII_TX1_N,
    SGMII_TX1_P,
    SPI_1_DO,
    USB_STP,
    // Inouts
    DQ,
    DQS,
    DQS_N,
    I2C_1_SCL,
    I2C_1_SDA,
    MAC_1_MDIO,
    QSPI_CLK,
    QSPI_DATA_0,
    QSPI_DATA_1,
    QSPI_DATA_2,
    QSPI_DATA_3,
    QSPI_SEL,
    RPi_GPIO12,
    RPi_GPIO13,
    RPi_GPIO16,
    RPi_GPIO17,
    RPi_GPIO19,
    RPi_GPIO20,
    RPi_GPIO21,
    RPi_GPIO22,
    RPi_GPIO23,
    RPi_GPIO24,
    RPi_GPIO25,
    RPi_GPIO26,
    RPi_GPIO27,
    SD_CMD_EMMC_CMD,
    SD_DATA0_EMMC_DATA0,
    SD_DATA1_EMMC_DATA1,
    SD_DATA2_EMMC_DATA2,
    SD_DATA3_EMMC_DATA3,
    SPI_1_CLK,
    SPI_1_SS0,
    USB_DATA0,
    USB_DATA1,
    USB_DATA2,
    USB_DATA3,
    USB_DATA4,
    USB_DATA5,
    USB_DATA6,
    USB_DATA7,
    mBUS_I2C_SCL,
    mBUS_I2C_SDA
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input         CAN_0_RXBUS_F2M;
input         CAN_1_RXBUS;
input         FIC_0_ACLK;
input         FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARREADY;
input         FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWREADY;
input  [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BID;
input  [1:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BRESP;
input         FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BVALID;
input  [63:0] FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RDATA;
input  [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RID;
input         FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RLAST;
input  [1:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RRESP;
input         FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RVALID;
input         FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WREADY;
input  [37:0] FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARADDR;
input  [1:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARBURST;
input  [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARCACHE;
input  [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARID;
input  [7:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLEN;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLOCK;
input  [2:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARPROT;
input  [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARQOS;
input  [2:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARSIZE;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARVALID;
input  [37:0] FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWADDR;
input  [1:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWBURST;
input  [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWCACHE;
input  [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWID;
input  [7:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLEN;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLOCK;
input  [2:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWPROT;
input  [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWQOS;
input  [2:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWSIZE;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWVALID;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BREADY;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RREADY;
input  [63:0] FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WDATA;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WLAST;
input  [7:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WSTRB;
input         FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WVALID;
input         FIC_1_ACLK;
input         FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARREADY;
input         FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWREADY;
input  [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BID;
input  [1:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BRESP;
input         FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BVALID;
input  [63:0] FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RDATA;
input  [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RID;
input         FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RLAST;
input  [1:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RRESP;
input         FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RVALID;
input         FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WREADY;
input  [37:0] FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARADDR;
input  [1:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARBURST;
input  [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARCACHE;
input  [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARID;
input  [7:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLEN;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLOCK;
input  [2:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARPROT;
input  [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARQOS;
input  [2:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARSIZE;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARVALID;
input  [37:0] FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWADDR;
input  [1:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWBURST;
input  [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWCACHE;
input  [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWID;
input  [7:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLEN;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLOCK;
input  [2:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWPROT;
input  [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWQOS;
input  [2:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWSIZE;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWVALID;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BREADY;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RREADY;
input  [63:0] FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WDATA;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WLAST;
input  [7:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WSTRB;
input         FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WVALID;
input         FIC_2_ACLK;
input  [37:0] FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARADDR;
input  [1:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARBURST;
input  [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARCACHE;
input  [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARID;
input  [7:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLEN;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLOCK;
input  [2:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARPROT;
input  [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARQOS;
input  [2:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARSIZE;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARVALID;
input  [37:0] FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWADDR;
input  [1:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWBURST;
input  [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWCACHE;
input  [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWID;
input  [7:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLEN;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLOCK;
input  [2:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWPROT;
input  [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWQOS;
input  [2:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWSIZE;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWVALID;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BREADY;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RREADY;
input  [63:0] FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WDATA;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WLAST;
input  [7:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WSTRB;
input         FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WVALID;
input  [31:0] FIC_3_APB_INITIATOR_FIC_3_APB_M_PRDATA;
input         FIC_3_APB_INITIATOR_FIC_3_APB_M_PREADY;
input         FIC_3_APB_INITIATOR_FIC_3_APB_M_PSLVERR;
input         FIC_3_PCLK;
input         GPIO_2_F2M_30;
input         GPIO_2_F2M_31;
input         MMUART_0_RXD_F2M;
input         MMUART_1_RXD_F2M;
input         MMUART_2_RXD_F2M;
input         MMUART_3_RXD_F2M;
input         MMUART_4_RXD_F2M;
input         MSS_INT_F2M_0;
input         MSS_INT_F2M_2;
input         MSS_INT_F2M_3;
input         MSS_RESET_N_F2M;
input         REFCLK;
input         REFCLK_N;
input         SD_CD_EMMC_STRB;
input         SD_WP_EMMC_RSTN;
input         SGMII_RX0_N;
input         SGMII_RX0_P;
input         SGMII_RX1_N;
input         SGMII_RX1_P;
input         SPI_1_DI;
input         USB_CLK;
input         USB_DIR;
input         USB_NXT;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [5:0]  CA;
output        CAN_0_TXBUS_M2F;
output        CAN_0_TX_EBL_M2F;
output        CAN_1_TXBUS;
output        CAN_1_TX_EBL_N;
output        CK;
output        CKE;
output        CK_N;
output        CS;
output [3:0]  DM;
output [37:0] FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARADDR;
output [1:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARBURST;
output [3:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARCACHE;
output [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARID;
output [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARLEN;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARLOCK;
output [2:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARPROT;
output [3:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARQOS;
output [2:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARSIZE;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARVALID;
output [37:0] FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWADDR;
output [1:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWBURST;
output [3:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWCACHE;
output [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWID;
output [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWLEN;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWLOCK;
output [2:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWPROT;
output [3:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWQOS;
output [2:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWSIZE;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWVALID;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BREADY;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RREADY;
output [63:0] FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WDATA;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WLAST;
output [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WSTRB;
output        FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WVALID;
output        FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARREADY;
output        FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWREADY;
output [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BID;
output [1:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BRESP;
output        FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BVALID;
output [63:0] FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RDATA;
output [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RID;
output        FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RLAST;
output [1:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RRESP;
output        FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RVALID;
output        FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WREADY;
output [37:0] FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARADDR;
output [1:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARBURST;
output [3:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARCACHE;
output [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARID;
output [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARLEN;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARLOCK;
output [2:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARPROT;
output [3:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARQOS;
output [2:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARSIZE;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARVALID;
output [37:0] FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWADDR;
output [1:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWBURST;
output [3:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWCACHE;
output [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWID;
output [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWLEN;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWLOCK;
output [2:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWPROT;
output [3:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWQOS;
output [2:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWSIZE;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWVALID;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BREADY;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RREADY;
output [63:0] FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WDATA;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WLAST;
output [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WSTRB;
output        FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WVALID;
output        FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARREADY;
output        FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWREADY;
output [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BID;
output [1:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BRESP;
output        FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BVALID;
output [63:0] FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RDATA;
output [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RID;
output        FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RLAST;
output [1:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RRESP;
output        FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RVALID;
output        FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WREADY;
output        FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARREADY;
output        FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWREADY;
output [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BID;
output [1:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BRESP;
output        FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BVALID;
output [63:0] FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RDATA;
output [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RID;
output        FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RLAST;
output [1:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RRESP;
output        FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RVALID;
output        FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WREADY;
output [28:0] FIC_3_APB_INITIATOR_FIC_3_APB_M_PADDR;
output        FIC_3_APB_INITIATOR_FIC_3_APB_M_PENABLE;
output        FIC_3_APB_INITIATOR_FIC_3_APB_M_PSEL;
output [31:0] FIC_3_APB_INITIATOR_FIC_3_APB_M_PWDATA;
output        FIC_3_APB_INITIATOR_FIC_3_APB_M_PWRITE;
output        GPIO_2_M2F_16;
output        GPIO_2_M2F_17;
output        GPIO_2_M2F_18;
output        GPIO_2_M2F_19;
output        GPIO_2_M2F_26;
output        GPIO_2_M2F_27;
output        GPIO_2_M2F_28;
output        MAC_1_MDC;
output        MMUART_0_TXD_M2F;
output        MMUART_1_TXD_M2F;
output        MMUART_2_TXD_M2F;
output        MMUART_3_TXD_M2F;
output        MMUART_4_TXD_M2F;
output        MSS_DLL_LOCKS;
output        MSS_RESET_N_M2F;
output        ODT;
output        RESET_N;
output        SD_CLK_EMMC_CLK;
output        SD_POW_EMMC_DATA4;
output        SD_VOLT_CMD_DIR_EMMC_DATA7;
output        SD_VOLT_DIR_0_EMMC_UNUSED;
output        SD_VOLT_DIR_1_3_EMMC_UNUSED;
output        SD_VOLT_EN_EMMC_DATA6;
output        SD_VOLT_SEL_EMMC_DATA5;
output        SGMII_TX0_N;
output        SGMII_TX0_P;
output        SGMII_TX1_N;
output        SGMII_TX1_P;
output        SPI_1_DO;
output        USB_STP;
//--------------------------------------------------------------------
// Inout
//--------------------------------------------------------------------
inout  [31:0] DQ;
inout  [3:0]  DQS;
inout  [3:0]  DQS_N;
inout         I2C_1_SCL;
inout         I2C_1_SDA;
inout         MAC_1_MDIO;
inout         QSPI_CLK;
inout         QSPI_DATA_0;
inout         QSPI_DATA_1;
inout         QSPI_DATA_2;
inout         QSPI_DATA_3;
inout         QSPI_SEL;
inout         RPi_GPIO12;
inout         RPi_GPIO13;
inout         RPi_GPIO16;
inout         RPi_GPIO17;
inout         RPi_GPIO19;
inout         RPi_GPIO20;
inout         RPi_GPIO21;
inout         RPi_GPIO22;
inout         RPi_GPIO23;
inout         RPi_GPIO24;
inout         RPi_GPIO25;
inout         RPi_GPIO26;
inout         RPi_GPIO27;
inout         SD_CMD_EMMC_CMD;
inout         SD_DATA0_EMMC_DATA0;
inout         SD_DATA1_EMMC_DATA1;
inout         SD_DATA2_EMMC_DATA2;
inout         SD_DATA3_EMMC_DATA3;
inout         SPI_1_CLK;
inout         SPI_1_SS0;
inout         USB_DATA0;
inout         USB_DATA1;
inout         USB_DATA2;
inout         USB_DATA3;
inout         USB_DATA4;
inout         USB_DATA5;
inout         USB_DATA6;
inout         USB_DATA7;
inout         mBUS_I2C_SCL;
inout         mBUS_I2C_SDA;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   [5:0]  CA_net_0;
wire          CAN_0_RXBUS_F2M;
wire          CAN_0_TX_EBL_M2F_net_0;
wire          CAN_0_TXBUS_M2F_net_0;
wire          CAN_1_RXBUS;
wire          CAN_1_TX_EBL_N_net_0;
wire          CAN_1_TXBUS_net_0;
wire          CK_net_0;
wire          CK_N_net_0;
wire          CKE_net_0;
wire          CS_net_0;
wire   [3:0]  DM_net_0;
wire   [31:0] DQ;
wire   [3:0]  DQS;
wire   [3:0]  DQS_N;
wire          FIC_0_ACLK;
wire   [37:0] FIC_0_AXI4_INITIATOR_ARADDR;
wire   [1:0]  FIC_0_AXI4_INITIATOR_ARBURST;
wire   [3:0]  FIC_0_AXI4_INITIATOR_ARCACHE;
wire   [7:0]  FIC_0_AXI4_INITIATOR_ARID;
wire   [7:0]  FIC_0_AXI4_INITIATOR_ARLEN;
wire          FIC_0_AXI4_INITIATOR_ARLOCK;
wire   [2:0]  FIC_0_AXI4_INITIATOR_ARPROT;
wire   [3:0]  FIC_0_AXI4_INITIATOR_ARQOS;
wire          FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARREADY;
wire   [2:0]  FIC_0_AXI4_INITIATOR_ARSIZE;
wire          FIC_0_AXI4_INITIATOR_ARVALID;
wire   [37:0] FIC_0_AXI4_INITIATOR_AWADDR;
wire   [1:0]  FIC_0_AXI4_INITIATOR_AWBURST;
wire   [3:0]  FIC_0_AXI4_INITIATOR_AWCACHE;
wire   [7:0]  FIC_0_AXI4_INITIATOR_AWID;
wire   [7:0]  FIC_0_AXI4_INITIATOR_AWLEN;
wire          FIC_0_AXI4_INITIATOR_AWLOCK;
wire   [2:0]  FIC_0_AXI4_INITIATOR_AWPROT;
wire   [3:0]  FIC_0_AXI4_INITIATOR_AWQOS;
wire          FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWREADY;
wire   [2:0]  FIC_0_AXI4_INITIATOR_AWSIZE;
wire          FIC_0_AXI4_INITIATOR_AWVALID;
wire   [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BID;
wire          FIC_0_AXI4_INITIATOR_BREADY;
wire   [1:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BRESP;
wire          FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BVALID;
wire   [63:0] FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RDATA;
wire   [7:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RID;
wire          FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RLAST;
wire          FIC_0_AXI4_INITIATOR_RREADY;
wire   [1:0]  FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RRESP;
wire          FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RVALID;
wire   [63:0] FIC_0_AXI4_INITIATOR_WDATA;
wire          FIC_0_AXI4_INITIATOR_WLAST;
wire          FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WREADY;
wire   [7:0]  FIC_0_AXI4_INITIATOR_WSTRB;
wire          FIC_0_AXI4_INITIATOR_WVALID;
wire   [37:0] FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARADDR;
wire   [1:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARBURST;
wire   [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARCACHE;
wire   [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARID;
wire   [7:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLEN;
wire          FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLOCK;
wire   [2:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARPROT;
wire   [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARQOS;
wire          FIC_0_AXI4_TARGET_ARREADY;
wire   [2:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARSIZE;
wire          FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARVALID;
wire   [37:0] FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWADDR;
wire   [1:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWBURST;
wire   [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWCACHE;
wire   [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWID;
wire   [7:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLEN;
wire          FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLOCK;
wire   [2:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWPROT;
wire   [3:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWQOS;
wire          FIC_0_AXI4_TARGET_AWREADY;
wire   [2:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWSIZE;
wire          FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWVALID;
wire   [3:0]  FIC_0_AXI4_TARGET_BID;
wire          FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BREADY;
wire   [1:0]  FIC_0_AXI4_TARGET_BRESP;
wire          FIC_0_AXI4_TARGET_BVALID;
wire   [63:0] FIC_0_AXI4_TARGET_RDATA;
wire   [3:0]  FIC_0_AXI4_TARGET_RID;
wire          FIC_0_AXI4_TARGET_RLAST;
wire          FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RREADY;
wire   [1:0]  FIC_0_AXI4_TARGET_RRESP;
wire          FIC_0_AXI4_TARGET_RVALID;
wire   [63:0] FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WDATA;
wire          FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WLAST;
wire          FIC_0_AXI4_TARGET_WREADY;
wire   [7:0]  FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WSTRB;
wire          FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WVALID;
wire          FIC_1_ACLK;
wire   [37:0] FIC_1_AXI4_INITIATOR_ARADDR;
wire   [1:0]  FIC_1_AXI4_INITIATOR_ARBURST;
wire   [3:0]  FIC_1_AXI4_INITIATOR_ARCACHE;
wire   [7:0]  FIC_1_AXI4_INITIATOR_ARID;
wire   [7:0]  FIC_1_AXI4_INITIATOR_ARLEN;
wire          FIC_1_AXI4_INITIATOR_ARLOCK;
wire   [2:0]  FIC_1_AXI4_INITIATOR_ARPROT;
wire   [3:0]  FIC_1_AXI4_INITIATOR_ARQOS;
wire          FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARREADY;
wire   [2:0]  FIC_1_AXI4_INITIATOR_ARSIZE;
wire          FIC_1_AXI4_INITIATOR_ARVALID;
wire   [37:0] FIC_1_AXI4_INITIATOR_AWADDR;
wire   [1:0]  FIC_1_AXI4_INITIATOR_AWBURST;
wire   [3:0]  FIC_1_AXI4_INITIATOR_AWCACHE;
wire   [7:0]  FIC_1_AXI4_INITIATOR_AWID;
wire   [7:0]  FIC_1_AXI4_INITIATOR_AWLEN;
wire          FIC_1_AXI4_INITIATOR_AWLOCK;
wire   [2:0]  FIC_1_AXI4_INITIATOR_AWPROT;
wire   [3:0]  FIC_1_AXI4_INITIATOR_AWQOS;
wire          FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWREADY;
wire   [2:0]  FIC_1_AXI4_INITIATOR_AWSIZE;
wire          FIC_1_AXI4_INITIATOR_AWVALID;
wire   [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BID;
wire          FIC_1_AXI4_INITIATOR_BREADY;
wire   [1:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BRESP;
wire          FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BVALID;
wire   [63:0] FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RDATA;
wire   [7:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RID;
wire          FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RLAST;
wire          FIC_1_AXI4_INITIATOR_RREADY;
wire   [1:0]  FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RRESP;
wire          FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RVALID;
wire   [63:0] FIC_1_AXI4_INITIATOR_WDATA;
wire          FIC_1_AXI4_INITIATOR_WLAST;
wire          FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WREADY;
wire   [7:0]  FIC_1_AXI4_INITIATOR_WSTRB;
wire          FIC_1_AXI4_INITIATOR_WVALID;
wire   [37:0] FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARADDR;
wire   [1:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARBURST;
wire   [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARCACHE;
wire   [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARID;
wire   [7:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLEN;
wire          FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLOCK;
wire   [2:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARPROT;
wire   [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARQOS;
wire          FIC_1_AXI4_TARGET_ARREADY;
wire   [2:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARSIZE;
wire          FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARVALID;
wire   [37:0] FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWADDR;
wire   [1:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWBURST;
wire   [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWCACHE;
wire   [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWID;
wire   [7:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLEN;
wire          FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLOCK;
wire   [2:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWPROT;
wire   [3:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWQOS;
wire          FIC_1_AXI4_TARGET_AWREADY;
wire   [2:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWSIZE;
wire          FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWVALID;
wire   [3:0]  FIC_1_AXI4_TARGET_BID;
wire          FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BREADY;
wire   [1:0]  FIC_1_AXI4_TARGET_BRESP;
wire          FIC_1_AXI4_TARGET_BVALID;
wire   [63:0] FIC_1_AXI4_TARGET_RDATA;
wire   [3:0]  FIC_1_AXI4_TARGET_RID;
wire          FIC_1_AXI4_TARGET_RLAST;
wire          FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RREADY;
wire   [1:0]  FIC_1_AXI4_TARGET_RRESP;
wire          FIC_1_AXI4_TARGET_RVALID;
wire   [63:0] FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WDATA;
wire          FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WLAST;
wire          FIC_1_AXI4_TARGET_WREADY;
wire   [7:0]  FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WSTRB;
wire          FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WVALID;
wire          FIC_2_ACLK;
wire   [37:0] FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARADDR;
wire   [1:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARBURST;
wire   [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARCACHE;
wire   [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARID;
wire   [7:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLEN;
wire          FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLOCK;
wire   [2:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARPROT;
wire   [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARQOS;
wire          FIC_2_AXI4_TARGET_ARREADY;
wire   [2:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARSIZE;
wire          FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARVALID;
wire   [37:0] FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWADDR;
wire   [1:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWBURST;
wire   [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWCACHE;
wire   [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWID;
wire   [7:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLEN;
wire          FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLOCK;
wire   [2:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWPROT;
wire   [3:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWQOS;
wire          FIC_2_AXI4_TARGET_AWREADY;
wire   [2:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWSIZE;
wire          FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWVALID;
wire   [3:0]  FIC_2_AXI4_TARGET_BID;
wire          FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BREADY;
wire   [1:0]  FIC_2_AXI4_TARGET_BRESP;
wire          FIC_2_AXI4_TARGET_BVALID;
wire   [63:0] FIC_2_AXI4_TARGET_RDATA;
wire   [3:0]  FIC_2_AXI4_TARGET_RID;
wire          FIC_2_AXI4_TARGET_RLAST;
wire          FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RREADY;
wire   [1:0]  FIC_2_AXI4_TARGET_RRESP;
wire          FIC_2_AXI4_TARGET_RVALID;
wire   [63:0] FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WDATA;
wire          FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WLAST;
wire          FIC_2_AXI4_TARGET_WREADY;
wire   [7:0]  FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WSTRB;
wire          FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WVALID;
wire   [28:0] FIC_3_APB_INITIATOR_PADDR;
wire          FIC_3_APB_INITIATOR_PENABLE;
wire   [31:0] FIC_3_APB_INITIATOR_FIC_3_APB_M_PRDATA;
wire          FIC_3_APB_INITIATOR_FIC_3_APB_M_PREADY;
wire          FIC_3_APB_INITIATOR_PSELx;
wire          FIC_3_APB_INITIATOR_FIC_3_APB_M_PSLVERR;
wire   [31:0] FIC_3_APB_INITIATOR_PWDATA;
wire          FIC_3_APB_INITIATOR_PWRITE;
wire          FIC_3_PCLK;
wire          GPIO_2_2_IO_Y;
wire          GPIO_2_3_IO_Y;
wire          GPIO_2_4_IO_Y;
wire          GPIO_2_5_IO_Y;
wire          GPIO_2_7_IO_Y;
wire          GPIO_2_8_IO_Y;
wire          GPIO_2_9_IO_Y;
wire          GPIO_2_10_IO_Y;
wire          GPIO_2_11_IO_Y;
wire          GPIO_2_12_IO_Y;
wire          GPIO_2_13_IO_Y;
wire          GPIO_2_14_IO_Y;
wire          GPIO_2_15_IO_Y;
wire          GPIO_2_F2M_30;
wire          GPIO_2_F2M_31;
wire          GPIO_2_M2F_16_net_0;
wire          GPIO_2_M2F_17_net_0;
wire          GPIO_2_M2F_18_net_0;
wire          GPIO_2_M2F_19_net_0;
wire          GPIO_2_M2F_26_net_0;
wire          GPIO_2_M2F_27_net_0;
wire          GPIO_2_M2F_28_net_0;
wire          I2C0_SCL_BIBUF_Y;
wire          I2C0_SDA_BIBUF_Y;
wire          I2C_1_SCL;
wire          I2C_1_SDA;
wire          ICICLE_MSS_FIC_0_DLL_LOCK_M2F;
wire          ICICLE_MSS_FIC_1_DLL_LOCK_M2F;
wire          ICICLE_MSS_FIC_2_DLL_LOCK_M2F;
wire          ICICLE_MSS_FIC_3_DLL_LOCK_M2F;
wire          ICICLE_MSS_GPIO_2_M2F_2;
wire          ICICLE_MSS_GPIO_2_M2F_3;
wire          ICICLE_MSS_GPIO_2_M2F_4;
wire          ICICLE_MSS_GPIO_2_M2F_5;
wire          ICICLE_MSS_GPIO_2_M2F_7;
wire          ICICLE_MSS_GPIO_2_M2F_8;
wire          ICICLE_MSS_GPIO_2_M2F_9;
wire          ICICLE_MSS_GPIO_2_M2F_10;
wire          ICICLE_MSS_GPIO_2_M2F_11;
wire          ICICLE_MSS_GPIO_2_M2F_12;
wire          ICICLE_MSS_GPIO_2_M2F_13;
wire          ICICLE_MSS_GPIO_2_M2F_14;
wire          ICICLE_MSS_GPIO_2_M2F_15;
wire          ICICLE_MSS_GPIO_2_OE_M2F_2;
wire          ICICLE_MSS_GPIO_2_OE_M2F_3;
wire          ICICLE_MSS_GPIO_2_OE_M2F_4;
wire          ICICLE_MSS_GPIO_2_OE_M2F_5;
wire          ICICLE_MSS_GPIO_2_OE_M2F_7;
wire          ICICLE_MSS_GPIO_2_OE_M2F_8;
wire          ICICLE_MSS_GPIO_2_OE_M2F_9;
wire          ICICLE_MSS_GPIO_2_OE_M2F_10;
wire          ICICLE_MSS_GPIO_2_OE_M2F_11;
wire          ICICLE_MSS_GPIO_2_OE_M2F_12;
wire          ICICLE_MSS_GPIO_2_OE_M2F_13;
wire          ICICLE_MSS_GPIO_2_OE_M2F_14;
wire          ICICLE_MSS_GPIO_2_OE_M2F_15;
wire          ICICLE_MSS_I2C_0_SCL_OE_M2F;
wire          ICICLE_MSS_I2C_0_SDA_OE_M2F;
wire          ICICLE_MSS_QSPI_CLK_M2F;
wire          ICICLE_MSS_QSPI_CLK_OE_M2F;
wire   [0:0]  ICICLE_MSS_QSPI_DATA_M2F0to0;
wire   [1:1]  ICICLE_MSS_QSPI_DATA_M2F1to1;
wire   [2:2]  ICICLE_MSS_QSPI_DATA_M2F2to2;
wire   [3:3]  ICICLE_MSS_QSPI_DATA_M2F3to3;
wire   [0:0]  ICICLE_MSS_QSPI_DATA_OE_M2F0to0;
wire   [1:1]  ICICLE_MSS_QSPI_DATA_OE_M2F1to1;
wire   [2:2]  ICICLE_MSS_QSPI_DATA_OE_M2F2to2;
wire   [3:3]  ICICLE_MSS_QSPI_DATA_OE_M2F3to3;
wire          ICICLE_MSS_QSPI_SEL_M2F;
wire          ICICLE_MSS_QSPI_SEL_OE_M2F;
wire          MAC_1_MDC_net_0;
wire          MAC_1_MDIO;
wire          mBUS_I2C_SCL;
wire          mBUS_I2C_SDA;
wire          MMUART_0_RXD_F2M;
wire          MMUART_0_TXD_M2F_net_0;
wire          MMUART_1_RXD_F2M;
wire          MMUART_1_TXD_M2F_net_0;
wire          MMUART_2_RXD_F2M;
wire          MMUART_2_TXD_M2F_net_0;
wire          MMUART_3_RXD_F2M;
wire          MMUART_3_TXD_M2F_net_0;
wire          MMUART_4_RXD_F2M;
wire          MMUART_4_TXD_M2F_net_0;
wire          MSS_DLL_LOCKS_net_0;
wire          MSS_INT_F2M_0;
wire          MSS_INT_F2M_2;
wire          MSS_INT_F2M_3;
wire          MSS_RESET_N_F2M;
wire          MSS_RESET_N_M2F_net_0;
wire          ODT_net_0;
wire          QSPI_CLK;
wire          QSPI_DATA_0;
wire          QSPI_DATA_0_BIBUF_Y;
wire          QSPI_DATA_1;
wire          QSPI_DATA_1_BIBUF_Y;
wire          QSPI_DATA_2;
wire          QSPI_DATA_2_BIBUF_Y;
wire          QSPI_DATA_3;
wire          QSPI_DATA_3_BIBUF_Y;
wire          QSPI_SEL;
wire          REFCLK;
wire          REFCLK_N;
wire          RESET_N_net_0;
wire          RPi_GPIO12;
wire          RPi_GPIO13;
wire          RPi_GPIO16;
wire          RPi_GPIO17;
wire          RPi_GPIO19;
wire          RPi_GPIO20;
wire          RPi_GPIO21;
wire          RPi_GPIO22;
wire          RPi_GPIO23;
wire          RPi_GPIO24;
wire          RPi_GPIO25;
wire          RPi_GPIO26;
wire          RPi_GPIO27;
wire          SD_CD_EMMC_STRB;
wire          SD_CLK_EMMC_CLK_net_0;
wire          SD_CMD_EMMC_CMD;
wire          SD_DATA0_EMMC_DATA0;
wire          SD_DATA1_EMMC_DATA1;
wire          SD_DATA2_EMMC_DATA2;
wire          SD_DATA3_EMMC_DATA3;
wire          SD_POW_EMMC_DATA4_net_0;
wire          SD_VOLT_CMD_DIR_EMMC_DATA7_net_0;
wire          SD_VOLT_DIR_0_EMMC_UNUSED_net_0;
wire          SD_VOLT_DIR_1_3_EMMC_UNUSED_net_0;
wire          SD_VOLT_EN_EMMC_DATA6_net_0;
wire          SD_VOLT_SEL_EMMC_DATA5_net_0;
wire          SD_WP_EMMC_RSTN;
wire          SGMII_RX0_N;
wire          SGMII_RX0_P;
wire          SGMII_RX1_N;
wire          SGMII_RX1_P;
wire          SGMII_TX0_N_net_0;
wire          SGMII_TX0_P_net_0;
wire          SGMII_TX1_N_net_0;
wire          SGMII_TX1_P_net_0;
wire          SPI_1_CLK;
wire          SPI_1_DI;
wire          SPI_1_DO_net_0;
wire          SPI_1_SS0;
wire          USB_CLK;
wire          USB_DATA0;
wire          USB_DATA1;
wire          USB_DATA2;
wire          USB_DATA3;
wire          USB_DATA4;
wire          USB_DATA5;
wire          USB_DATA6;
wire          USB_DATA7;
wire          USB_DIR;
wire          USB_NXT;
wire          USB_STP_net_0;
wire          CAN_0_TXBUS_M2F_net_1;
wire          CAN_0_TX_EBL_M2F_net_1;
wire          CAN_1_TXBUS_net_1;
wire          CAN_1_TX_EBL_N_net_1;
wire          CKE_net_1;
wire          CK_N_net_1;
wire          CK_net_1;
wire          CS_net_1;
wire          FIC_0_AXI4_INITIATOR_ARLOCK_net_0;
wire          FIC_0_AXI4_INITIATOR_ARVALID_net_0;
wire          FIC_0_AXI4_INITIATOR_AWLOCK_net_0;
wire          FIC_0_AXI4_INITIATOR_AWVALID_net_0;
wire          FIC_0_AXI4_INITIATOR_BREADY_net_0;
wire          FIC_0_AXI4_INITIATOR_RREADY_net_0;
wire          FIC_0_AXI4_INITIATOR_WLAST_net_0;
wire          FIC_0_AXI4_INITIATOR_WVALID_net_0;
wire          FIC_0_AXI4_TARGET_ARREADY_net_0;
wire          FIC_0_AXI4_TARGET_AWREADY_net_0;
wire          FIC_0_AXI4_TARGET_BVALID_net_0;
wire          FIC_0_AXI4_TARGET_RLAST_net_0;
wire          FIC_0_AXI4_TARGET_RVALID_net_0;
wire          FIC_0_AXI4_TARGET_WREADY_net_0;
wire          FIC_1_AXI4_INITIATOR_ARLOCK_net_0;
wire          FIC_1_AXI4_INITIATOR_ARVALID_net_0;
wire          FIC_1_AXI4_INITIATOR_AWLOCK_net_0;
wire          FIC_1_AXI4_INITIATOR_AWVALID_net_0;
wire          FIC_1_AXI4_INITIATOR_BREADY_net_0;
wire          FIC_1_AXI4_INITIATOR_RREADY_net_0;
wire          FIC_1_AXI4_INITIATOR_WLAST_net_0;
wire          FIC_1_AXI4_INITIATOR_WVALID_net_0;
wire          FIC_1_AXI4_TARGET_ARREADY_net_0;
wire          FIC_1_AXI4_TARGET_AWREADY_net_0;
wire          FIC_1_AXI4_TARGET_BVALID_net_0;
wire          FIC_1_AXI4_TARGET_RLAST_net_0;
wire          FIC_1_AXI4_TARGET_RVALID_net_0;
wire          FIC_1_AXI4_TARGET_WREADY_net_0;
wire          FIC_2_AXI4_TARGET_ARREADY_net_0;
wire          FIC_2_AXI4_TARGET_AWREADY_net_0;
wire          FIC_2_AXI4_TARGET_BVALID_net_0;
wire          FIC_2_AXI4_TARGET_RLAST_net_0;
wire          FIC_2_AXI4_TARGET_RVALID_net_0;
wire          FIC_2_AXI4_TARGET_WREADY_net_0;
wire          FIC_3_APB_INITIATOR_PENABLE_net_0;
wire          FIC_3_APB_INITIATOR_PSELx_net_0;
wire          FIC_3_APB_INITIATOR_PWRITE_net_0;
wire          GPIO_2_M2F_16_net_1;
wire          GPIO_2_M2F_17_net_1;
wire          GPIO_2_M2F_18_net_1;
wire          GPIO_2_M2F_19_net_1;
wire          GPIO_2_M2F_26_net_1;
wire          GPIO_2_M2F_27_net_1;
wire          GPIO_2_M2F_28_net_1;
wire          MAC_1_MDC_net_1;
wire          MMUART_0_TXD_M2F_net_1;
wire          MMUART_1_TXD_M2F_net_1;
wire          MMUART_2_TXD_M2F_net_1;
wire          MMUART_3_TXD_M2F_net_1;
wire          MMUART_4_TXD_M2F_net_1;
wire          MSS_DLL_LOCKS_net_1;
wire          MSS_RESET_N_M2F_net_1;
wire          ODT_net_1;
wire          RESET_N_net_1;
wire          SD_CLK_EMMC_CLK_net_1;
wire          SD_POW_EMMC_DATA4_net_1;
wire          SD_VOLT_CMD_DIR_EMMC_DATA7_net_1;
wire          SD_VOLT_DIR_0_EMMC_UNUSED_net_1;
wire          SD_VOLT_DIR_1_3_EMMC_UNUSED_net_1;
wire          SD_VOLT_EN_EMMC_DATA6_net_1;
wire          SD_VOLT_SEL_EMMC_DATA5_net_1;
wire          SGMII_TX0_N_net_1;
wire          SGMII_TX0_P_net_1;
wire          SGMII_TX1_N_net_1;
wire          SGMII_TX1_P_net_1;
wire          SPI_1_DO_net_1;
wire          USB_STP_net_1;
wire   [5:0]  CA_net_1;
wire   [3:0]  DM_net_1;
wire   [37:0] FIC_0_AXI4_INITIATOR_ARADDR_net_0;
wire   [1:0]  FIC_0_AXI4_INITIATOR_ARBURST_net_0;
wire   [3:0]  FIC_0_AXI4_INITIATOR_ARCACHE_net_0;
wire   [7:0]  FIC_0_AXI4_INITIATOR_ARID_net_0;
wire   [7:0]  FIC_0_AXI4_INITIATOR_ARLEN_net_0;
wire   [2:0]  FIC_0_AXI4_INITIATOR_ARPROT_net_0;
wire   [3:0]  FIC_0_AXI4_INITIATOR_ARQOS_net_0;
wire   [2:0]  FIC_0_AXI4_INITIATOR_ARSIZE_net_0;
wire   [37:0] FIC_0_AXI4_INITIATOR_AWADDR_net_0;
wire   [1:0]  FIC_0_AXI4_INITIATOR_AWBURST_net_0;
wire   [3:0]  FIC_0_AXI4_INITIATOR_AWCACHE_net_0;
wire   [7:0]  FIC_0_AXI4_INITIATOR_AWID_net_0;
wire   [7:0]  FIC_0_AXI4_INITIATOR_AWLEN_net_0;
wire   [2:0]  FIC_0_AXI4_INITIATOR_AWPROT_net_0;
wire   [3:0]  FIC_0_AXI4_INITIATOR_AWQOS_net_0;
wire   [2:0]  FIC_0_AXI4_INITIATOR_AWSIZE_net_0;
wire   [63:0] FIC_0_AXI4_INITIATOR_WDATA_net_0;
wire   [7:0]  FIC_0_AXI4_INITIATOR_WSTRB_net_0;
wire   [3:0]  FIC_0_AXI4_TARGET_BID_net_0;
wire   [1:0]  FIC_0_AXI4_TARGET_BRESP_net_0;
wire   [63:0] FIC_0_AXI4_TARGET_RDATA_net_0;
wire   [3:0]  FIC_0_AXI4_TARGET_RID_net_0;
wire   [1:0]  FIC_0_AXI4_TARGET_RRESP_net_0;
wire   [37:0] FIC_1_AXI4_INITIATOR_ARADDR_net_0;
wire   [1:0]  FIC_1_AXI4_INITIATOR_ARBURST_net_0;
wire   [3:0]  FIC_1_AXI4_INITIATOR_ARCACHE_net_0;
wire   [7:0]  FIC_1_AXI4_INITIATOR_ARID_net_0;
wire   [7:0]  FIC_1_AXI4_INITIATOR_ARLEN_net_0;
wire   [2:0]  FIC_1_AXI4_INITIATOR_ARPROT_net_0;
wire   [3:0]  FIC_1_AXI4_INITIATOR_ARQOS_net_0;
wire   [2:0]  FIC_1_AXI4_INITIATOR_ARSIZE_net_0;
wire   [37:0] FIC_1_AXI4_INITIATOR_AWADDR_net_0;
wire   [1:0]  FIC_1_AXI4_INITIATOR_AWBURST_net_0;
wire   [3:0]  FIC_1_AXI4_INITIATOR_AWCACHE_net_0;
wire   [7:0]  FIC_1_AXI4_INITIATOR_AWID_net_0;
wire   [7:0]  FIC_1_AXI4_INITIATOR_AWLEN_net_0;
wire   [2:0]  FIC_1_AXI4_INITIATOR_AWPROT_net_0;
wire   [3:0]  FIC_1_AXI4_INITIATOR_AWQOS_net_0;
wire   [2:0]  FIC_1_AXI4_INITIATOR_AWSIZE_net_0;
wire   [63:0] FIC_1_AXI4_INITIATOR_WDATA_net_0;
wire   [7:0]  FIC_1_AXI4_INITIATOR_WSTRB_net_0;
wire   [3:0]  FIC_1_AXI4_TARGET_BID_net_0;
wire   [1:0]  FIC_1_AXI4_TARGET_BRESP_net_0;
wire   [63:0] FIC_1_AXI4_TARGET_RDATA_net_0;
wire   [3:0]  FIC_1_AXI4_TARGET_RID_net_0;
wire   [1:0]  FIC_1_AXI4_TARGET_RRESP_net_0;
wire   [3:0]  FIC_2_AXI4_TARGET_BID_net_0;
wire   [1:0]  FIC_2_AXI4_TARGET_BRESP_net_0;
wire   [63:0] FIC_2_AXI4_TARGET_RDATA_net_0;
wire   [3:0]  FIC_2_AXI4_TARGET_RID_net_0;
wire   [1:0]  FIC_2_AXI4_TARGET_RRESP_net_0;
wire   [28:0] FIC_3_APB_INITIATOR_PADDR_net_0;
wire   [31:0] FIC_3_APB_INITIATOR_PWDATA_net_0;
wire   [3:0]  QSPI_DATA_F2M_net_0;
wire   [63:0] MSS_INT_F2M_net_0;
wire   [3:0]  QSPI_DATA_M2F_net_0;
wire   [3:0]  QSPI_DATA_OE_M2F_net_0;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire          GND_net;
wire   [63:4] MSS_INT_F2M_const_net_0;
//--------------------------------------------------------------------
// Inverted Nets
//--------------------------------------------------------------------
wire          CAN_0_TX_EBL_M2F_OUT_PRE_INV0_0;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign GND_net                 = 1'b0;
assign MSS_INT_F2M_const_net_0 = 60'h000000000000000;
//--------------------------------------------------------------------
// Inversions
//--------------------------------------------------------------------
assign CAN_0_TX_EBL_M2F_net_0 = ~ CAN_0_TX_EBL_M2F_OUT_PRE_INV0_0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign CAN_0_TXBUS_M2F_net_1                          = CAN_0_TXBUS_M2F_net_0;
assign CAN_0_TXBUS_M2F                                = CAN_0_TXBUS_M2F_net_1;
assign CAN_0_TX_EBL_M2F_net_1                         = CAN_0_TX_EBL_M2F_net_0;
assign CAN_0_TX_EBL_M2F                               = CAN_0_TX_EBL_M2F_net_1;
assign CAN_1_TXBUS_net_1                              = CAN_1_TXBUS_net_0;
assign CAN_1_TXBUS                                    = CAN_1_TXBUS_net_1;
assign CAN_1_TX_EBL_N_net_1                           = CAN_1_TX_EBL_N_net_0;
assign CAN_1_TX_EBL_N                                 = CAN_1_TX_EBL_N_net_1;
assign CKE_net_1                                      = CKE_net_0;
assign CKE                                            = CKE_net_1;
assign CK_N_net_1                                     = CK_N_net_0;
assign CK_N                                           = CK_N_net_1;
assign CK_net_1                                       = CK_net_0;
assign CK                                             = CK_net_1;
assign CS_net_1                                       = CS_net_0;
assign CS                                             = CS_net_1;
assign FIC_0_AXI4_INITIATOR_ARLOCK_net_0              = FIC_0_AXI4_INITIATOR_ARLOCK;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARLOCK       = FIC_0_AXI4_INITIATOR_ARLOCK_net_0;
assign FIC_0_AXI4_INITIATOR_ARVALID_net_0             = FIC_0_AXI4_INITIATOR_ARVALID;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARVALID      = FIC_0_AXI4_INITIATOR_ARVALID_net_0;
assign FIC_0_AXI4_INITIATOR_AWLOCK_net_0              = FIC_0_AXI4_INITIATOR_AWLOCK;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWLOCK       = FIC_0_AXI4_INITIATOR_AWLOCK_net_0;
assign FIC_0_AXI4_INITIATOR_AWVALID_net_0             = FIC_0_AXI4_INITIATOR_AWVALID;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWVALID      = FIC_0_AXI4_INITIATOR_AWVALID_net_0;
assign FIC_0_AXI4_INITIATOR_BREADY_net_0              = FIC_0_AXI4_INITIATOR_BREADY;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BREADY       = FIC_0_AXI4_INITIATOR_BREADY_net_0;
assign FIC_0_AXI4_INITIATOR_RREADY_net_0              = FIC_0_AXI4_INITIATOR_RREADY;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RREADY       = FIC_0_AXI4_INITIATOR_RREADY_net_0;
assign FIC_0_AXI4_INITIATOR_WLAST_net_0               = FIC_0_AXI4_INITIATOR_WLAST;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WLAST        = FIC_0_AXI4_INITIATOR_WLAST_net_0;
assign FIC_0_AXI4_INITIATOR_WVALID_net_0              = FIC_0_AXI4_INITIATOR_WVALID;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WVALID       = FIC_0_AXI4_INITIATOR_WVALID_net_0;
assign FIC_0_AXI4_TARGET_ARREADY_net_0                = FIC_0_AXI4_TARGET_ARREADY;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARREADY         = FIC_0_AXI4_TARGET_ARREADY_net_0;
assign FIC_0_AXI4_TARGET_AWREADY_net_0                = FIC_0_AXI4_TARGET_AWREADY;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWREADY         = FIC_0_AXI4_TARGET_AWREADY_net_0;
assign FIC_0_AXI4_TARGET_BVALID_net_0                 = FIC_0_AXI4_TARGET_BVALID;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BVALID          = FIC_0_AXI4_TARGET_BVALID_net_0;
assign FIC_0_AXI4_TARGET_RLAST_net_0                  = FIC_0_AXI4_TARGET_RLAST;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RLAST           = FIC_0_AXI4_TARGET_RLAST_net_0;
assign FIC_0_AXI4_TARGET_RVALID_net_0                 = FIC_0_AXI4_TARGET_RVALID;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RVALID          = FIC_0_AXI4_TARGET_RVALID_net_0;
assign FIC_0_AXI4_TARGET_WREADY_net_0                 = FIC_0_AXI4_TARGET_WREADY;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WREADY          = FIC_0_AXI4_TARGET_WREADY_net_0;
assign FIC_1_AXI4_INITIATOR_ARLOCK_net_0              = FIC_1_AXI4_INITIATOR_ARLOCK;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARLOCK       = FIC_1_AXI4_INITIATOR_ARLOCK_net_0;
assign FIC_1_AXI4_INITIATOR_ARVALID_net_0             = FIC_1_AXI4_INITIATOR_ARVALID;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARVALID      = FIC_1_AXI4_INITIATOR_ARVALID_net_0;
assign FIC_1_AXI4_INITIATOR_AWLOCK_net_0              = FIC_1_AXI4_INITIATOR_AWLOCK;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWLOCK       = FIC_1_AXI4_INITIATOR_AWLOCK_net_0;
assign FIC_1_AXI4_INITIATOR_AWVALID_net_0             = FIC_1_AXI4_INITIATOR_AWVALID;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWVALID      = FIC_1_AXI4_INITIATOR_AWVALID_net_0;
assign FIC_1_AXI4_INITIATOR_BREADY_net_0              = FIC_1_AXI4_INITIATOR_BREADY;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BREADY       = FIC_1_AXI4_INITIATOR_BREADY_net_0;
assign FIC_1_AXI4_INITIATOR_RREADY_net_0              = FIC_1_AXI4_INITIATOR_RREADY;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RREADY       = FIC_1_AXI4_INITIATOR_RREADY_net_0;
assign FIC_1_AXI4_INITIATOR_WLAST_net_0               = FIC_1_AXI4_INITIATOR_WLAST;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WLAST        = FIC_1_AXI4_INITIATOR_WLAST_net_0;
assign FIC_1_AXI4_INITIATOR_WVALID_net_0              = FIC_1_AXI4_INITIATOR_WVALID;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WVALID       = FIC_1_AXI4_INITIATOR_WVALID_net_0;
assign FIC_1_AXI4_TARGET_ARREADY_net_0                = FIC_1_AXI4_TARGET_ARREADY;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARREADY         = FIC_1_AXI4_TARGET_ARREADY_net_0;
assign FIC_1_AXI4_TARGET_AWREADY_net_0                = FIC_1_AXI4_TARGET_AWREADY;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWREADY         = FIC_1_AXI4_TARGET_AWREADY_net_0;
assign FIC_1_AXI4_TARGET_BVALID_net_0                 = FIC_1_AXI4_TARGET_BVALID;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BVALID          = FIC_1_AXI4_TARGET_BVALID_net_0;
assign FIC_1_AXI4_TARGET_RLAST_net_0                  = FIC_1_AXI4_TARGET_RLAST;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RLAST           = FIC_1_AXI4_TARGET_RLAST_net_0;
assign FIC_1_AXI4_TARGET_RVALID_net_0                 = FIC_1_AXI4_TARGET_RVALID;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RVALID          = FIC_1_AXI4_TARGET_RVALID_net_0;
assign FIC_1_AXI4_TARGET_WREADY_net_0                 = FIC_1_AXI4_TARGET_WREADY;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WREADY          = FIC_1_AXI4_TARGET_WREADY_net_0;
assign FIC_2_AXI4_TARGET_ARREADY_net_0                = FIC_2_AXI4_TARGET_ARREADY;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARREADY         = FIC_2_AXI4_TARGET_ARREADY_net_0;
assign FIC_2_AXI4_TARGET_AWREADY_net_0                = FIC_2_AXI4_TARGET_AWREADY;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWREADY         = FIC_2_AXI4_TARGET_AWREADY_net_0;
assign FIC_2_AXI4_TARGET_BVALID_net_0                 = FIC_2_AXI4_TARGET_BVALID;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BVALID          = FIC_2_AXI4_TARGET_BVALID_net_0;
assign FIC_2_AXI4_TARGET_RLAST_net_0                  = FIC_2_AXI4_TARGET_RLAST;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RLAST           = FIC_2_AXI4_TARGET_RLAST_net_0;
assign FIC_2_AXI4_TARGET_RVALID_net_0                 = FIC_2_AXI4_TARGET_RVALID;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RVALID          = FIC_2_AXI4_TARGET_RVALID_net_0;
assign FIC_2_AXI4_TARGET_WREADY_net_0                 = FIC_2_AXI4_TARGET_WREADY;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WREADY          = FIC_2_AXI4_TARGET_WREADY_net_0;
assign FIC_3_APB_INITIATOR_PENABLE_net_0              = FIC_3_APB_INITIATOR_PENABLE;
assign FIC_3_APB_INITIATOR_FIC_3_APB_M_PENABLE        = FIC_3_APB_INITIATOR_PENABLE_net_0;
assign FIC_3_APB_INITIATOR_PSELx_net_0                = FIC_3_APB_INITIATOR_PSELx;
assign FIC_3_APB_INITIATOR_FIC_3_APB_M_PSEL           = FIC_3_APB_INITIATOR_PSELx_net_0;
assign FIC_3_APB_INITIATOR_PWRITE_net_0               = FIC_3_APB_INITIATOR_PWRITE;
assign FIC_3_APB_INITIATOR_FIC_3_APB_M_PWRITE         = FIC_3_APB_INITIATOR_PWRITE_net_0;
assign GPIO_2_M2F_16_net_1                            = GPIO_2_M2F_16_net_0;
assign GPIO_2_M2F_16                                  = GPIO_2_M2F_16_net_1;
assign GPIO_2_M2F_17_net_1                            = GPIO_2_M2F_17_net_0;
assign GPIO_2_M2F_17                                  = GPIO_2_M2F_17_net_1;
assign GPIO_2_M2F_18_net_1                            = GPIO_2_M2F_18_net_0;
assign GPIO_2_M2F_18                                  = GPIO_2_M2F_18_net_1;
assign GPIO_2_M2F_19_net_1                            = GPIO_2_M2F_19_net_0;
assign GPIO_2_M2F_19                                  = GPIO_2_M2F_19_net_1;
assign GPIO_2_M2F_26_net_1                            = GPIO_2_M2F_26_net_0;
assign GPIO_2_M2F_26                                  = GPIO_2_M2F_26_net_1;
assign GPIO_2_M2F_27_net_1                            = GPIO_2_M2F_27_net_0;
assign GPIO_2_M2F_27                                  = GPIO_2_M2F_27_net_1;
assign GPIO_2_M2F_28_net_1                            = GPIO_2_M2F_28_net_0;
assign GPIO_2_M2F_28                                  = GPIO_2_M2F_28_net_1;
assign MAC_1_MDC_net_1                                = MAC_1_MDC_net_0;
assign MAC_1_MDC                                      = MAC_1_MDC_net_1;
assign MMUART_0_TXD_M2F_net_1                         = MMUART_0_TXD_M2F_net_0;
assign MMUART_0_TXD_M2F                               = MMUART_0_TXD_M2F_net_1;
assign MMUART_1_TXD_M2F_net_1                         = MMUART_1_TXD_M2F_net_0;
assign MMUART_1_TXD_M2F                               = MMUART_1_TXD_M2F_net_1;
assign MMUART_2_TXD_M2F_net_1                         = MMUART_2_TXD_M2F_net_0;
assign MMUART_2_TXD_M2F                               = MMUART_2_TXD_M2F_net_1;
assign MMUART_3_TXD_M2F_net_1                         = MMUART_3_TXD_M2F_net_0;
assign MMUART_3_TXD_M2F                               = MMUART_3_TXD_M2F_net_1;
assign MMUART_4_TXD_M2F_net_1                         = MMUART_4_TXD_M2F_net_0;
assign MMUART_4_TXD_M2F                               = MMUART_4_TXD_M2F_net_1;
assign MSS_DLL_LOCKS_net_1                            = MSS_DLL_LOCKS_net_0;
assign MSS_DLL_LOCKS                                  = MSS_DLL_LOCKS_net_1;
assign MSS_RESET_N_M2F_net_1                          = MSS_RESET_N_M2F_net_0;
assign MSS_RESET_N_M2F                                = MSS_RESET_N_M2F_net_1;
assign ODT_net_1                                      = ODT_net_0;
assign ODT                                            = ODT_net_1;
assign RESET_N_net_1                                  = RESET_N_net_0;
assign RESET_N                                        = RESET_N_net_1;
assign SD_CLK_EMMC_CLK_net_1                          = SD_CLK_EMMC_CLK_net_0;
assign SD_CLK_EMMC_CLK                                = SD_CLK_EMMC_CLK_net_1;
assign SD_POW_EMMC_DATA4_net_1                        = SD_POW_EMMC_DATA4_net_0;
assign SD_POW_EMMC_DATA4                              = SD_POW_EMMC_DATA4_net_1;
assign SD_VOLT_CMD_DIR_EMMC_DATA7_net_1               = SD_VOLT_CMD_DIR_EMMC_DATA7_net_0;
assign SD_VOLT_CMD_DIR_EMMC_DATA7                     = SD_VOLT_CMD_DIR_EMMC_DATA7_net_1;
assign SD_VOLT_DIR_0_EMMC_UNUSED_net_1                = SD_VOLT_DIR_0_EMMC_UNUSED_net_0;
assign SD_VOLT_DIR_0_EMMC_UNUSED                      = SD_VOLT_DIR_0_EMMC_UNUSED_net_1;
assign SD_VOLT_DIR_1_3_EMMC_UNUSED_net_1              = SD_VOLT_DIR_1_3_EMMC_UNUSED_net_0;
assign SD_VOLT_DIR_1_3_EMMC_UNUSED                    = SD_VOLT_DIR_1_3_EMMC_UNUSED_net_1;
assign SD_VOLT_EN_EMMC_DATA6_net_1                    = SD_VOLT_EN_EMMC_DATA6_net_0;
assign SD_VOLT_EN_EMMC_DATA6                          = SD_VOLT_EN_EMMC_DATA6_net_1;
assign SD_VOLT_SEL_EMMC_DATA5_net_1                   = SD_VOLT_SEL_EMMC_DATA5_net_0;
assign SD_VOLT_SEL_EMMC_DATA5                         = SD_VOLT_SEL_EMMC_DATA5_net_1;
assign SGMII_TX0_N_net_1                              = SGMII_TX0_N_net_0;
assign SGMII_TX0_N                                    = SGMII_TX0_N_net_1;
assign SGMII_TX0_P_net_1                              = SGMII_TX0_P_net_0;
assign SGMII_TX0_P                                    = SGMII_TX0_P_net_1;
assign SGMII_TX1_N_net_1                              = SGMII_TX1_N_net_0;
assign SGMII_TX1_N                                    = SGMII_TX1_N_net_1;
assign SGMII_TX1_P_net_1                              = SGMII_TX1_P_net_0;
assign SGMII_TX1_P                                    = SGMII_TX1_P_net_1;
assign SPI_1_DO_net_1                                 = SPI_1_DO_net_0;
assign SPI_1_DO                                       = SPI_1_DO_net_1;
assign USB_STP_net_1                                  = USB_STP_net_0;
assign USB_STP                                        = USB_STP_net_1;
assign CA_net_1                                       = CA_net_0;
assign CA[5:0]                                        = CA_net_1;
assign DM_net_1                                       = DM_net_0;
assign DM[3:0]                                        = DM_net_1;
assign FIC_0_AXI4_INITIATOR_ARADDR_net_0              = FIC_0_AXI4_INITIATOR_ARADDR;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARADDR[37:0] = FIC_0_AXI4_INITIATOR_ARADDR_net_0;
assign FIC_0_AXI4_INITIATOR_ARBURST_net_0             = FIC_0_AXI4_INITIATOR_ARBURST;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARBURST[1:0] = FIC_0_AXI4_INITIATOR_ARBURST_net_0;
assign FIC_0_AXI4_INITIATOR_ARCACHE_net_0             = FIC_0_AXI4_INITIATOR_ARCACHE;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARCACHE[3:0] = FIC_0_AXI4_INITIATOR_ARCACHE_net_0;
assign FIC_0_AXI4_INITIATOR_ARID_net_0                = FIC_0_AXI4_INITIATOR_ARID;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARID[7:0]    = FIC_0_AXI4_INITIATOR_ARID_net_0;
assign FIC_0_AXI4_INITIATOR_ARLEN_net_0               = FIC_0_AXI4_INITIATOR_ARLEN;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARLEN[7:0]   = FIC_0_AXI4_INITIATOR_ARLEN_net_0;
assign FIC_0_AXI4_INITIATOR_ARPROT_net_0              = FIC_0_AXI4_INITIATOR_ARPROT;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARPROT[2:0]  = FIC_0_AXI4_INITIATOR_ARPROT_net_0;
assign FIC_0_AXI4_INITIATOR_ARQOS_net_0               = FIC_0_AXI4_INITIATOR_ARQOS;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARQOS[3:0]   = FIC_0_AXI4_INITIATOR_ARQOS_net_0;
assign FIC_0_AXI4_INITIATOR_ARSIZE_net_0              = FIC_0_AXI4_INITIATOR_ARSIZE;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARSIZE[2:0]  = FIC_0_AXI4_INITIATOR_ARSIZE_net_0;
assign FIC_0_AXI4_INITIATOR_AWADDR_net_0              = FIC_0_AXI4_INITIATOR_AWADDR;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWADDR[37:0] = FIC_0_AXI4_INITIATOR_AWADDR_net_0;
assign FIC_0_AXI4_INITIATOR_AWBURST_net_0             = FIC_0_AXI4_INITIATOR_AWBURST;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWBURST[1:0] = FIC_0_AXI4_INITIATOR_AWBURST_net_0;
assign FIC_0_AXI4_INITIATOR_AWCACHE_net_0             = FIC_0_AXI4_INITIATOR_AWCACHE;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWCACHE[3:0] = FIC_0_AXI4_INITIATOR_AWCACHE_net_0;
assign FIC_0_AXI4_INITIATOR_AWID_net_0                = FIC_0_AXI4_INITIATOR_AWID;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWID[7:0]    = FIC_0_AXI4_INITIATOR_AWID_net_0;
assign FIC_0_AXI4_INITIATOR_AWLEN_net_0               = FIC_0_AXI4_INITIATOR_AWLEN;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWLEN[7:0]   = FIC_0_AXI4_INITIATOR_AWLEN_net_0;
assign FIC_0_AXI4_INITIATOR_AWPROT_net_0              = FIC_0_AXI4_INITIATOR_AWPROT;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWPROT[2:0]  = FIC_0_AXI4_INITIATOR_AWPROT_net_0;
assign FIC_0_AXI4_INITIATOR_AWQOS_net_0               = FIC_0_AXI4_INITIATOR_AWQOS;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWQOS[3:0]   = FIC_0_AXI4_INITIATOR_AWQOS_net_0;
assign FIC_0_AXI4_INITIATOR_AWSIZE_net_0              = FIC_0_AXI4_INITIATOR_AWSIZE;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWSIZE[2:0]  = FIC_0_AXI4_INITIATOR_AWSIZE_net_0;
assign FIC_0_AXI4_INITIATOR_WDATA_net_0               = FIC_0_AXI4_INITIATOR_WDATA;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WDATA[63:0]  = FIC_0_AXI4_INITIATOR_WDATA_net_0;
assign FIC_0_AXI4_INITIATOR_WSTRB_net_0               = FIC_0_AXI4_INITIATOR_WSTRB;
assign FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WSTRB[7:0]   = FIC_0_AXI4_INITIATOR_WSTRB_net_0;
assign FIC_0_AXI4_TARGET_BID_net_0                    = FIC_0_AXI4_TARGET_BID;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BID[3:0]        = FIC_0_AXI4_TARGET_BID_net_0;
assign FIC_0_AXI4_TARGET_BRESP_net_0                  = FIC_0_AXI4_TARGET_BRESP;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BRESP[1:0]      = FIC_0_AXI4_TARGET_BRESP_net_0;
assign FIC_0_AXI4_TARGET_RDATA_net_0                  = FIC_0_AXI4_TARGET_RDATA;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RDATA[63:0]     = FIC_0_AXI4_TARGET_RDATA_net_0;
assign FIC_0_AXI4_TARGET_RID_net_0                    = FIC_0_AXI4_TARGET_RID;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RID[3:0]        = FIC_0_AXI4_TARGET_RID_net_0;
assign FIC_0_AXI4_TARGET_RRESP_net_0                  = FIC_0_AXI4_TARGET_RRESP;
assign FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RRESP[1:0]      = FIC_0_AXI4_TARGET_RRESP_net_0;
assign FIC_1_AXI4_INITIATOR_ARADDR_net_0              = FIC_1_AXI4_INITIATOR_ARADDR;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARADDR[37:0] = FIC_1_AXI4_INITIATOR_ARADDR_net_0;
assign FIC_1_AXI4_INITIATOR_ARBURST_net_0             = FIC_1_AXI4_INITIATOR_ARBURST;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARBURST[1:0] = FIC_1_AXI4_INITIATOR_ARBURST_net_0;
assign FIC_1_AXI4_INITIATOR_ARCACHE_net_0             = FIC_1_AXI4_INITIATOR_ARCACHE;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARCACHE[3:0] = FIC_1_AXI4_INITIATOR_ARCACHE_net_0;
assign FIC_1_AXI4_INITIATOR_ARID_net_0                = FIC_1_AXI4_INITIATOR_ARID;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARID[7:0]    = FIC_1_AXI4_INITIATOR_ARID_net_0;
assign FIC_1_AXI4_INITIATOR_ARLEN_net_0               = FIC_1_AXI4_INITIATOR_ARLEN;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARLEN[7:0]   = FIC_1_AXI4_INITIATOR_ARLEN_net_0;
assign FIC_1_AXI4_INITIATOR_ARPROT_net_0              = FIC_1_AXI4_INITIATOR_ARPROT;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARPROT[2:0]  = FIC_1_AXI4_INITIATOR_ARPROT_net_0;
assign FIC_1_AXI4_INITIATOR_ARQOS_net_0               = FIC_1_AXI4_INITIATOR_ARQOS;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARQOS[3:0]   = FIC_1_AXI4_INITIATOR_ARQOS_net_0;
assign FIC_1_AXI4_INITIATOR_ARSIZE_net_0              = FIC_1_AXI4_INITIATOR_ARSIZE;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARSIZE[2:0]  = FIC_1_AXI4_INITIATOR_ARSIZE_net_0;
assign FIC_1_AXI4_INITIATOR_AWADDR_net_0              = FIC_1_AXI4_INITIATOR_AWADDR;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWADDR[37:0] = FIC_1_AXI4_INITIATOR_AWADDR_net_0;
assign FIC_1_AXI4_INITIATOR_AWBURST_net_0             = FIC_1_AXI4_INITIATOR_AWBURST;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWBURST[1:0] = FIC_1_AXI4_INITIATOR_AWBURST_net_0;
assign FIC_1_AXI4_INITIATOR_AWCACHE_net_0             = FIC_1_AXI4_INITIATOR_AWCACHE;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWCACHE[3:0] = FIC_1_AXI4_INITIATOR_AWCACHE_net_0;
assign FIC_1_AXI4_INITIATOR_AWID_net_0                = FIC_1_AXI4_INITIATOR_AWID;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWID[7:0]    = FIC_1_AXI4_INITIATOR_AWID_net_0;
assign FIC_1_AXI4_INITIATOR_AWLEN_net_0               = FIC_1_AXI4_INITIATOR_AWLEN;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWLEN[7:0]   = FIC_1_AXI4_INITIATOR_AWLEN_net_0;
assign FIC_1_AXI4_INITIATOR_AWPROT_net_0              = FIC_1_AXI4_INITIATOR_AWPROT;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWPROT[2:0]  = FIC_1_AXI4_INITIATOR_AWPROT_net_0;
assign FIC_1_AXI4_INITIATOR_AWQOS_net_0               = FIC_1_AXI4_INITIATOR_AWQOS;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWQOS[3:0]   = FIC_1_AXI4_INITIATOR_AWQOS_net_0;
assign FIC_1_AXI4_INITIATOR_AWSIZE_net_0              = FIC_1_AXI4_INITIATOR_AWSIZE;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWSIZE[2:0]  = FIC_1_AXI4_INITIATOR_AWSIZE_net_0;
assign FIC_1_AXI4_INITIATOR_WDATA_net_0               = FIC_1_AXI4_INITIATOR_WDATA;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WDATA[63:0]  = FIC_1_AXI4_INITIATOR_WDATA_net_0;
assign FIC_1_AXI4_INITIATOR_WSTRB_net_0               = FIC_1_AXI4_INITIATOR_WSTRB;
assign FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WSTRB[7:0]   = FIC_1_AXI4_INITIATOR_WSTRB_net_0;
assign FIC_1_AXI4_TARGET_BID_net_0                    = FIC_1_AXI4_TARGET_BID;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BID[3:0]        = FIC_1_AXI4_TARGET_BID_net_0;
assign FIC_1_AXI4_TARGET_BRESP_net_0                  = FIC_1_AXI4_TARGET_BRESP;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BRESP[1:0]      = FIC_1_AXI4_TARGET_BRESP_net_0;
assign FIC_1_AXI4_TARGET_RDATA_net_0                  = FIC_1_AXI4_TARGET_RDATA;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RDATA[63:0]     = FIC_1_AXI4_TARGET_RDATA_net_0;
assign FIC_1_AXI4_TARGET_RID_net_0                    = FIC_1_AXI4_TARGET_RID;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RID[3:0]        = FIC_1_AXI4_TARGET_RID_net_0;
assign FIC_1_AXI4_TARGET_RRESP_net_0                  = FIC_1_AXI4_TARGET_RRESP;
assign FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RRESP[1:0]      = FIC_1_AXI4_TARGET_RRESP_net_0;
assign FIC_2_AXI4_TARGET_BID_net_0                    = FIC_2_AXI4_TARGET_BID;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BID[3:0]        = FIC_2_AXI4_TARGET_BID_net_0;
assign FIC_2_AXI4_TARGET_BRESP_net_0                  = FIC_2_AXI4_TARGET_BRESP;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BRESP[1:0]      = FIC_2_AXI4_TARGET_BRESP_net_0;
assign FIC_2_AXI4_TARGET_RDATA_net_0                  = FIC_2_AXI4_TARGET_RDATA;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RDATA[63:0]     = FIC_2_AXI4_TARGET_RDATA_net_0;
assign FIC_2_AXI4_TARGET_RID_net_0                    = FIC_2_AXI4_TARGET_RID;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RID[3:0]        = FIC_2_AXI4_TARGET_RID_net_0;
assign FIC_2_AXI4_TARGET_RRESP_net_0                  = FIC_2_AXI4_TARGET_RRESP;
assign FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RRESP[1:0]      = FIC_2_AXI4_TARGET_RRESP_net_0;
assign FIC_3_APB_INITIATOR_PADDR_net_0                = FIC_3_APB_INITIATOR_PADDR;
assign FIC_3_APB_INITIATOR_FIC_3_APB_M_PADDR[28:0]    = FIC_3_APB_INITIATOR_PADDR_net_0;
assign FIC_3_APB_INITIATOR_PWDATA_net_0               = FIC_3_APB_INITIATOR_PWDATA;
assign FIC_3_APB_INITIATOR_FIC_3_APB_M_PWDATA[31:0]   = FIC_3_APB_INITIATOR_PWDATA_net_0;
//--------------------------------------------------------------------
// Slices assignments
//--------------------------------------------------------------------
assign ICICLE_MSS_QSPI_DATA_M2F0to0[0]    = QSPI_DATA_M2F_net_0[0:0];
assign ICICLE_MSS_QSPI_DATA_M2F1to1[1]    = QSPI_DATA_M2F_net_0[1:1];
assign ICICLE_MSS_QSPI_DATA_M2F2to2[2]    = QSPI_DATA_M2F_net_0[2:2];
assign ICICLE_MSS_QSPI_DATA_M2F3to3[3]    = QSPI_DATA_M2F_net_0[3:3];
assign ICICLE_MSS_QSPI_DATA_OE_M2F0to0[0] = QSPI_DATA_OE_M2F_net_0[0:0];
assign ICICLE_MSS_QSPI_DATA_OE_M2F1to1[1] = QSPI_DATA_OE_M2F_net_0[1:1];
assign ICICLE_MSS_QSPI_DATA_OE_M2F2to2[2] = QSPI_DATA_OE_M2F_net_0[2:2];
assign ICICLE_MSS_QSPI_DATA_OE_M2F3to3[3] = QSPI_DATA_OE_M2F_net_0[3:3];
//--------------------------------------------------------------------
// Concatenation assignments
//--------------------------------------------------------------------
assign QSPI_DATA_F2M_net_0 = { QSPI_DATA_3_BIBUF_Y , QSPI_DATA_2_BIBUF_Y , QSPI_DATA_1_BIBUF_Y , QSPI_DATA_0_BIBUF_Y };
assign MSS_INT_F2M_net_0   = { 60'h000000000000000 , MSS_INT_F2M_3 , MSS_INT_F2M_2 , 1'b0 , MSS_INT_F2M_0 };
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------AND4
AND4 AND4_MSS_DLL_LOCKS(
        // Inputs
        .A ( ICICLE_MSS_FIC_0_DLL_LOCK_M2F ),
        .B ( ICICLE_MSS_FIC_3_DLL_LOCK_M2F ),
        .C ( ICICLE_MSS_FIC_2_DLL_LOCK_M2F ),
        .D ( ICICLE_MSS_FIC_1_DLL_LOCK_M2F ),
        // Outputs
        .Y ( MSS_DLL_LOCKS_net_0 ) 
        );

//--------BIBUF
BIBUF GPIO_2_2_IO(
        // Inputs
        .D   ( ICICLE_MSS_GPIO_2_M2F_2 ),
        .E   ( ICICLE_MSS_GPIO_2_OE_M2F_2 ),
        // Outputs
        .Y   ( GPIO_2_2_IO_Y ),
        // Inouts
        .PAD ( RPi_GPIO12 ) 
        );

//--------BIBUF
BIBUF GPIO_2_3_IO(
        // Inputs
        .D   ( ICICLE_MSS_GPIO_2_M2F_3 ),
        .E   ( ICICLE_MSS_GPIO_2_OE_M2F_3 ),
        // Outputs
        .Y   ( GPIO_2_3_IO_Y ),
        // Inouts
        .PAD ( RPi_GPIO13 ) 
        );

//--------BIBUF
BIBUF GPIO_2_4_IO(
        // Inputs
        .D   ( ICICLE_MSS_GPIO_2_M2F_4 ),
        .E   ( ICICLE_MSS_GPIO_2_OE_M2F_4 ),
        // Outputs
        .Y   ( GPIO_2_4_IO_Y ),
        // Inouts
        .PAD ( RPi_GPIO16 ) 
        );

//--------BIBUF
BIBUF GPIO_2_5_IO(
        // Inputs
        .D   ( ICICLE_MSS_GPIO_2_M2F_5 ),
        .E   ( ICICLE_MSS_GPIO_2_OE_M2F_5 ),
        // Outputs
        .Y   ( GPIO_2_5_IO_Y ),
        // Inouts
        .PAD ( RPi_GPIO17 ) 
        );

//--------BIBUF
BIBUF GPIO_2_7_IO(
        // Inputs
        .D   ( ICICLE_MSS_GPIO_2_M2F_7 ),
        .E   ( ICICLE_MSS_GPIO_2_OE_M2F_7 ),
        // Outputs
        .Y   ( GPIO_2_7_IO_Y ),
        // Inouts
        .PAD ( RPi_GPIO19 ) 
        );

//--------BIBUF
BIBUF GPIO_2_8_IO(
        // Inputs
        .D   ( ICICLE_MSS_GPIO_2_M2F_8 ),
        .E   ( ICICLE_MSS_GPIO_2_OE_M2F_8 ),
        // Outputs
        .Y   ( GPIO_2_8_IO_Y ),
        // Inouts
        .PAD ( RPi_GPIO20 ) 
        );

//--------BIBUF
BIBUF GPIO_2_9_IO(
        // Inputs
        .D   ( ICICLE_MSS_GPIO_2_M2F_9 ),
        .E   ( ICICLE_MSS_GPIO_2_OE_M2F_9 ),
        // Outputs
        .Y   ( GPIO_2_9_IO_Y ),
        // Inouts
        .PAD ( RPi_GPIO21 ) 
        );

//--------BIBUF
BIBUF GPIO_2_10_IO(
        // Inputs
        .D   ( ICICLE_MSS_GPIO_2_M2F_10 ),
        .E   ( ICICLE_MSS_GPIO_2_OE_M2F_10 ),
        // Outputs
        .Y   ( GPIO_2_10_IO_Y ),
        // Inouts
        .PAD ( RPi_GPIO22 ) 
        );

//--------BIBUF
BIBUF GPIO_2_11_IO(
        // Inputs
        .D   ( ICICLE_MSS_GPIO_2_M2F_11 ),
        .E   ( ICICLE_MSS_GPIO_2_OE_M2F_11 ),
        // Outputs
        .Y   ( GPIO_2_11_IO_Y ),
        // Inouts
        .PAD ( RPi_GPIO23 ) 
        );

//--------BIBUF
BIBUF GPIO_2_12_IO(
        // Inputs
        .D   ( ICICLE_MSS_GPIO_2_M2F_12 ),
        .E   ( ICICLE_MSS_GPIO_2_OE_M2F_12 ),
        // Outputs
        .Y   ( GPIO_2_12_IO_Y ),
        // Inouts
        .PAD ( RPi_GPIO24 ) 
        );

//--------BIBUF
BIBUF GPIO_2_13_IO(
        // Inputs
        .D   ( ICICLE_MSS_GPIO_2_M2F_13 ),
        .E   ( ICICLE_MSS_GPIO_2_OE_M2F_13 ),
        // Outputs
        .Y   ( GPIO_2_13_IO_Y ),
        // Inouts
        .PAD ( RPi_GPIO25 ) 
        );

//--------BIBUF
BIBUF GPIO_2_14_IO(
        // Inputs
        .D   ( ICICLE_MSS_GPIO_2_M2F_14 ),
        .E   ( ICICLE_MSS_GPIO_2_OE_M2F_14 ),
        // Outputs
        .Y   ( GPIO_2_14_IO_Y ),
        // Inouts
        .PAD ( RPi_GPIO26 ) 
        );

//--------BIBUF
BIBUF GPIO_2_15_IO(
        // Inputs
        .D   ( ICICLE_MSS_GPIO_2_M2F_15 ),
        .E   ( ICICLE_MSS_GPIO_2_OE_M2F_15 ),
        // Outputs
        .Y   ( GPIO_2_15_IO_Y ),
        // Inouts
        .PAD ( RPi_GPIO27 ) 
        );

//--------BIBUF
BIBUF I2C0_SCL_BIBUF(
        // Inputs
        .D   ( GND_net ),
        .E   ( ICICLE_MSS_I2C_0_SCL_OE_M2F ),
        // Outputs
        .Y   ( I2C0_SCL_BIBUF_Y ),
        // Inouts
        .PAD ( mBUS_I2C_SCL ) 
        );

//--------BIBUF
BIBUF I2C0_SDA_BIBUF(
        // Inputs
        .D   ( GND_net ),
        .E   ( ICICLE_MSS_I2C_0_SDA_OE_M2F ),
        // Outputs
        .Y   ( I2C0_SDA_BIBUF_Y ),
        // Inouts
        .PAD ( mBUS_I2C_SDA ) 
        );

//--------ICICLE_MSS
ICICLE_MSS ICICLE_MSS_inst_0(
        // Inputs
        .FIC_0_ACLK                   ( FIC_0_ACLK ),
        .FIC_0_AXI4_M_AWREADY         ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_AWREADY ),
        .FIC_0_AXI4_M_WREADY          ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_WREADY ),
        .FIC_0_AXI4_M_BVALID          ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BVALID ),
        .FIC_0_AXI4_M_ARREADY         ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_ARREADY ),
        .FIC_0_AXI4_M_RLAST           ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RLAST ),
        .FIC_0_AXI4_M_RVALID          ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RVALID ),
        .FIC_0_AXI4_S_AWLOCK          ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLOCK ),
        .FIC_0_AXI4_S_AWVALID         ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWVALID ),
        .FIC_0_AXI4_S_WLAST           ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WLAST ),
        .FIC_0_AXI4_S_WVALID          ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WVALID ),
        .FIC_0_AXI4_S_BREADY          ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_BREADY ),
        .FIC_0_AXI4_S_ARLOCK          ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLOCK ),
        .FIC_0_AXI4_S_ARVALID         ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARVALID ),
        .FIC_0_AXI4_S_RREADY          ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_RREADY ),
        .FIC_1_ACLK                   ( FIC_1_ACLK ),
        .FIC_1_AXI4_M_AWREADY         ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_AWREADY ),
        .FIC_1_AXI4_M_WREADY          ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_WREADY ),
        .FIC_1_AXI4_M_BVALID          ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BVALID ),
        .FIC_1_AXI4_M_ARREADY         ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_ARREADY ),
        .FIC_1_AXI4_M_RLAST           ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RLAST ),
        .FIC_1_AXI4_M_RVALID          ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RVALID ),
        .FIC_1_AXI4_S_AWLOCK          ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLOCK ),
        .FIC_1_AXI4_S_AWVALID         ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWVALID ),
        .FIC_1_AXI4_S_WLAST           ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WLAST ),
        .FIC_1_AXI4_S_WVALID          ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WVALID ),
        .FIC_1_AXI4_S_BREADY          ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_BREADY ),
        .FIC_1_AXI4_S_ARLOCK          ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLOCK ),
        .FIC_1_AXI4_S_ARVALID         ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARVALID ),
        .FIC_1_AXI4_S_RREADY          ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_RREADY ),
        .FIC_2_ACLK                   ( FIC_2_ACLK ),
        .FIC_2_AXI4_S_AWLOCK          ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLOCK ),
        .FIC_2_AXI4_S_AWVALID         ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWVALID ),
        .FIC_2_AXI4_S_WLAST           ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WLAST ),
        .FIC_2_AXI4_S_WVALID          ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WVALID ),
        .FIC_2_AXI4_S_BREADY          ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_BREADY ),
        .FIC_2_AXI4_S_ARLOCK          ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLOCK ),
        .FIC_2_AXI4_S_ARVALID         ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARVALID ),
        .FIC_2_AXI4_S_RREADY          ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_RREADY ),
        .FIC_3_PCLK                   ( FIC_3_PCLK ),
        .FIC_3_APB_M_PREADY           ( FIC_3_APB_INITIATOR_FIC_3_APB_M_PREADY ),
        .FIC_3_APB_M_PSLVERR          ( FIC_3_APB_INITIATOR_FIC_3_APB_M_PSLVERR ),
        .MMUART_0_RXD_F2M             ( MMUART_0_RXD_F2M ),
        .MMUART_1_RXD_F2M             ( MMUART_1_RXD_F2M ),
        .MMUART_2_RXD_F2M             ( MMUART_2_RXD_F2M ),
        .MMUART_3_RXD_F2M             ( MMUART_3_RXD_F2M ),
        .MMUART_4_RXD_F2M             ( MMUART_4_RXD_F2M ),
        .CAN_0_RXBUS_F2M              ( CAN_0_RXBUS_F2M ),
        .SPI_0_SS_F2M                 ( GND_net ),
        .SPI_0_DI_F2M                 ( GND_net ),
        .SPI_0_CLK_F2M                ( GND_net ),
        .I2C_0_SCL_F2M                ( I2C0_SCL_BIBUF_Y ),
        .I2C_0_SDA_F2M                ( I2C0_SDA_BIBUF_Y ),
        .GPIO_2_F2M_31                ( GPIO_2_F2M_31 ),
        .GPIO_2_F2M_30                ( GPIO_2_F2M_30 ),
        .GPIO_2_F2M_15                ( GPIO_2_15_IO_Y ),
        .GPIO_2_F2M_14                ( GPIO_2_14_IO_Y ),
        .GPIO_2_F2M_13                ( GPIO_2_13_IO_Y ),
        .GPIO_2_F2M_12                ( GPIO_2_12_IO_Y ),
        .GPIO_2_F2M_11                ( GPIO_2_11_IO_Y ),
        .GPIO_2_F2M_10                ( GPIO_2_10_IO_Y ),
        .GPIO_2_F2M_9                 ( GPIO_2_9_IO_Y ),
        .GPIO_2_F2M_8                 ( GPIO_2_8_IO_Y ),
        .GPIO_2_F2M_7                 ( GPIO_2_7_IO_Y ),
        .GPIO_2_F2M_6                 ( GND_net ),
        .GPIO_2_F2M_5                 ( GPIO_2_5_IO_Y ),
        .GPIO_2_F2M_4                 ( GPIO_2_4_IO_Y ),
        .GPIO_2_F2M_3                 ( GPIO_2_3_IO_Y ),
        .GPIO_2_F2M_2                 ( GPIO_2_2_IO_Y ),
        .GPIO_2_F2M_1                 ( GND_net ),
        .GPIO_2_F2M_0                 ( GND_net ),
        .MSS_RESET_N_F2M              ( MSS_RESET_N_F2M ),
        .CAN_1_RXBUS                  ( CAN_1_RXBUS ),
        .USB_CLK                      ( USB_CLK ),
        .USB_DIR                      ( USB_DIR ),
        .USB_NXT                      ( USB_NXT ),
        .SPI_1_DI                     ( SPI_1_DI ),
        .SD_CD_EMMC_STRB              ( SD_CD_EMMC_STRB ),
        .SD_WP_EMMC_RSTN              ( SD_WP_EMMC_RSTN ),
        .SGMII_RX1_P                  ( SGMII_RX1_P ),
        .SGMII_RX1_N                  ( SGMII_RX1_N ),
        .SGMII_RX0_P                  ( SGMII_RX0_P ),
        .SGMII_RX0_N                  ( SGMII_RX0_N ),
        .REFCLK                       ( REFCLK ),
        .REFCLK_N                     ( REFCLK_N ),
        .FIC_0_AXI4_M_BID             ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BID ),
        .FIC_0_AXI4_M_BRESP           ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_BRESP ),
        .FIC_0_AXI4_M_RID             ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RID ),
        .FIC_0_AXI4_M_RDATA           ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RDATA ),
        .FIC_0_AXI4_M_RRESP           ( FIC_0_AXI4_INITIATOR_FIC_0_AXI4_M_RRESP ),
        .FIC_0_AXI4_S_AWID            ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWID ),
        .FIC_0_AXI4_S_AWADDR          ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWADDR ),
        .FIC_0_AXI4_S_AWLEN           ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWLEN ),
        .FIC_0_AXI4_S_AWSIZE          ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWSIZE ),
        .FIC_0_AXI4_S_AWBURST         ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWBURST ),
        .FIC_0_AXI4_S_AWQOS           ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWQOS ),
        .FIC_0_AXI4_S_AWCACHE         ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWCACHE ),
        .FIC_0_AXI4_S_AWPROT          ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_AWPROT ),
        .FIC_0_AXI4_S_WDATA           ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WDATA ),
        .FIC_0_AXI4_S_WSTRB           ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_WSTRB ),
        .FIC_0_AXI4_S_ARID            ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARID ),
        .FIC_0_AXI4_S_ARADDR          ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARADDR ),
        .FIC_0_AXI4_S_ARLEN           ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARLEN ),
        .FIC_0_AXI4_S_ARSIZE          ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARSIZE ),
        .FIC_0_AXI4_S_ARBURST         ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARBURST ),
        .FIC_0_AXI4_S_ARQOS           ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARQOS ),
        .FIC_0_AXI4_S_ARCACHE         ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARCACHE ),
        .FIC_0_AXI4_S_ARPROT          ( FIC_0_AXI4_TARGET_FIC_0_AXI4_S_ARPROT ),
        .FIC_1_AXI4_M_BID             ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BID ),
        .FIC_1_AXI4_M_BRESP           ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_BRESP ),
        .FIC_1_AXI4_M_RID             ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RID ),
        .FIC_1_AXI4_M_RDATA           ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RDATA ),
        .FIC_1_AXI4_M_RRESP           ( FIC_1_AXI4_INITIATOR_FIC_1_AXI4_M_RRESP ),
        .FIC_1_AXI4_S_AWID            ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWID ),
        .FIC_1_AXI4_S_AWADDR          ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWADDR ),
        .FIC_1_AXI4_S_AWLEN           ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWLEN ),
        .FIC_1_AXI4_S_AWSIZE          ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWSIZE ),
        .FIC_1_AXI4_S_AWBURST         ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWBURST ),
        .FIC_1_AXI4_S_AWCACHE         ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWCACHE ),
        .FIC_1_AXI4_S_AWQOS           ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWQOS ),
        .FIC_1_AXI4_S_AWPROT          ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_AWPROT ),
        .FIC_1_AXI4_S_WDATA           ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WDATA ),
        .FIC_1_AXI4_S_WSTRB           ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_WSTRB ),
        .FIC_1_AXI4_S_ARID            ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARID ),
        .FIC_1_AXI4_S_ARADDR          ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARADDR ),
        .FIC_1_AXI4_S_ARLEN           ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARLEN ),
        .FIC_1_AXI4_S_ARSIZE          ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARSIZE ),
        .FIC_1_AXI4_S_ARBURST         ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARBURST ),
        .FIC_1_AXI4_S_ARQOS           ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARQOS ),
        .FIC_1_AXI4_S_ARCACHE         ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARCACHE ),
        .FIC_1_AXI4_S_ARPROT          ( FIC_1_AXI4_TARGET_FIC_1_AXI4_S_ARPROT ),
        .FIC_2_AXI4_S_AWID            ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWID ),
        .FIC_2_AXI4_S_AWADDR          ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWADDR ),
        .FIC_2_AXI4_S_AWLEN           ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWLEN ),
        .FIC_2_AXI4_S_AWSIZE          ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWSIZE ),
        .FIC_2_AXI4_S_AWBURST         ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWBURST ),
        .FIC_2_AXI4_S_AWCACHE         ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWCACHE ),
        .FIC_2_AXI4_S_AWQOS           ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWQOS ),
        .FIC_2_AXI4_S_AWPROT          ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_AWPROT ),
        .FIC_2_AXI4_S_WDATA           ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WDATA ),
        .FIC_2_AXI4_S_WSTRB           ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_WSTRB ),
        .FIC_2_AXI4_S_ARID            ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARID ),
        .FIC_2_AXI4_S_ARADDR          ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARADDR ),
        .FIC_2_AXI4_S_ARLEN           ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARLEN ),
        .FIC_2_AXI4_S_ARSIZE          ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARSIZE ),
        .FIC_2_AXI4_S_ARBURST         ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARBURST ),
        .FIC_2_AXI4_S_ARCACHE         ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARCACHE ),
        .FIC_2_AXI4_S_ARQOS           ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARQOS ),
        .FIC_2_AXI4_S_ARPROT          ( FIC_2_AXI4_TARGET_FIC_2_AXI4_S_ARPROT ),
        .FIC_3_APB_M_PRDATA           ( FIC_3_APB_INITIATOR_FIC_3_APB_M_PRDATA ),
        .QSPI_DATA_F2M                ( QSPI_DATA_F2M_net_0 ),
        .MSS_INT_F2M                  ( MSS_INT_F2M_net_0 ),
        // Outputs
        .FIC_0_DLL_LOCK_M2F           ( ICICLE_MSS_FIC_0_DLL_LOCK_M2F ),
        .FIC_1_DLL_LOCK_M2F           ( ICICLE_MSS_FIC_1_DLL_LOCK_M2F ),
        .FIC_2_DLL_LOCK_M2F           ( ICICLE_MSS_FIC_2_DLL_LOCK_M2F ),
        .FIC_3_DLL_LOCK_M2F           ( ICICLE_MSS_FIC_3_DLL_LOCK_M2F ),
        .FIC_0_AXI4_M_AWLOCK          ( FIC_0_AXI4_INITIATOR_AWLOCK ),
        .FIC_0_AXI4_M_AWVALID         ( FIC_0_AXI4_INITIATOR_AWVALID ),
        .FIC_0_AXI4_M_WLAST           ( FIC_0_AXI4_INITIATOR_WLAST ),
        .FIC_0_AXI4_M_WVALID          ( FIC_0_AXI4_INITIATOR_WVALID ),
        .FIC_0_AXI4_M_BREADY          ( FIC_0_AXI4_INITIATOR_BREADY ),
        .FIC_0_AXI4_M_ARLOCK          ( FIC_0_AXI4_INITIATOR_ARLOCK ),
        .FIC_0_AXI4_M_ARVALID         ( FIC_0_AXI4_INITIATOR_ARVALID ),
        .FIC_0_AXI4_M_RREADY          ( FIC_0_AXI4_INITIATOR_RREADY ),
        .FIC_0_AXI4_S_AWREADY         ( FIC_0_AXI4_TARGET_AWREADY ),
        .FIC_0_AXI4_S_WREADY          ( FIC_0_AXI4_TARGET_WREADY ),
        .FIC_0_AXI4_S_BVALID          ( FIC_0_AXI4_TARGET_BVALID ),
        .FIC_0_AXI4_S_ARREADY         ( FIC_0_AXI4_TARGET_ARREADY ),
        .FIC_0_AXI4_S_RLAST           ( FIC_0_AXI4_TARGET_RLAST ),
        .FIC_0_AXI4_S_RVALID          ( FIC_0_AXI4_TARGET_RVALID ),
        .FIC_1_AXI4_M_AWLOCK          ( FIC_1_AXI4_INITIATOR_AWLOCK ),
        .FIC_1_AXI4_M_AWVALID         ( FIC_1_AXI4_INITIATOR_AWVALID ),
        .FIC_1_AXI4_M_WLAST           ( FIC_1_AXI4_INITIATOR_WLAST ),
        .FIC_1_AXI4_M_WVALID          ( FIC_1_AXI4_INITIATOR_WVALID ),
        .FIC_1_AXI4_M_BREADY          ( FIC_1_AXI4_INITIATOR_BREADY ),
        .FIC_1_AXI4_M_ARLOCK          ( FIC_1_AXI4_INITIATOR_ARLOCK ),
        .FIC_1_AXI4_M_ARVALID         ( FIC_1_AXI4_INITIATOR_ARVALID ),
        .FIC_1_AXI4_M_RREADY          ( FIC_1_AXI4_INITIATOR_RREADY ),
        .FIC_1_AXI4_S_AWREADY         ( FIC_1_AXI4_TARGET_AWREADY ),
        .FIC_1_AXI4_S_WREADY          ( FIC_1_AXI4_TARGET_WREADY ),
        .FIC_1_AXI4_S_BVALID          ( FIC_1_AXI4_TARGET_BVALID ),
        .FIC_1_AXI4_S_ARREADY         ( FIC_1_AXI4_TARGET_ARREADY ),
        .FIC_1_AXI4_S_RLAST           ( FIC_1_AXI4_TARGET_RLAST ),
        .FIC_1_AXI4_S_RVALID          ( FIC_1_AXI4_TARGET_RVALID ),
        .FIC_2_AXI4_S_AWREADY         ( FIC_2_AXI4_TARGET_AWREADY ),
        .FIC_2_AXI4_S_WREADY          ( FIC_2_AXI4_TARGET_WREADY ),
        .FIC_2_AXI4_S_BVALID          ( FIC_2_AXI4_TARGET_BVALID ),
        .FIC_2_AXI4_S_ARREADY         ( FIC_2_AXI4_TARGET_ARREADY ),
        .FIC_2_AXI4_S_RLAST           ( FIC_2_AXI4_TARGET_RLAST ),
        .FIC_2_AXI4_S_RVALID          ( FIC_2_AXI4_TARGET_RVALID ),
        .FIC_3_APB_M_PSEL             ( FIC_3_APB_INITIATOR_PSELx ),
        .FIC_3_APB_M_PWRITE           ( FIC_3_APB_INITIATOR_PWRITE ),
        .FIC_3_APB_M_PENABLE          ( FIC_3_APB_INITIATOR_PENABLE ),
        .MMUART_0_TXD_M2F             ( MMUART_0_TXD_M2F_net_0 ),
        .MMUART_0_TXD_OE_M2F          (  ),
        .MMUART_1_TXD_M2F             ( MMUART_1_TXD_M2F_net_0 ),
        .MMUART_1_TXD_OE_M2F          (  ),
        .MMUART_2_TXD_M2F             ( MMUART_2_TXD_M2F_net_0 ),
        .MMUART_3_TXD_M2F             ( MMUART_3_TXD_M2F_net_0 ),
        .MMUART_4_TXD_M2F             ( MMUART_4_TXD_M2F_net_0 ),
        .CAN_0_TX_EBL_M2F             ( CAN_0_TX_EBL_M2F_OUT_PRE_INV0_0 ),
        .CAN_0_TXBUS_M2F              ( CAN_0_TXBUS_M2F_net_0 ),
        .QSPI_SEL_M2F                 ( ICICLE_MSS_QSPI_SEL_M2F ),
        .QSPI_SEL_OE_M2F              ( ICICLE_MSS_QSPI_SEL_OE_M2F ),
        .QSPI_CLK_M2F                 ( ICICLE_MSS_QSPI_CLK_M2F ),
        .QSPI_CLK_OE_M2F              ( ICICLE_MSS_QSPI_CLK_OE_M2F ),
        .SPI_0_SS1_M2F                (  ),
        .SPI_0_SS1_OE_M2F             (  ),
        .SPI_0_DO_M2F                 (  ),
        .SPI_0_DO_OE_M2F              (  ),
        .SPI_0_CLK_M2F                (  ),
        .SPI_0_CLK_OE_M2F             (  ),
        .I2C_0_SCL_OE_M2F             ( ICICLE_MSS_I2C_0_SCL_OE_M2F ),
        .I2C_0_SDA_OE_M2F             ( ICICLE_MSS_I2C_0_SDA_OE_M2F ),
        .GPIO_2_M2F_28                ( GPIO_2_M2F_28_net_0 ),
        .GPIO_2_M2F_27                ( GPIO_2_M2F_27_net_0 ),
        .GPIO_2_M2F_26                ( GPIO_2_M2F_26_net_0 ),
        .GPIO_2_M2F_19                ( GPIO_2_M2F_19_net_0 ),
        .GPIO_2_M2F_18                ( GPIO_2_M2F_18_net_0 ),
        .GPIO_2_M2F_17                ( GPIO_2_M2F_17_net_0 ),
        .GPIO_2_M2F_16                ( GPIO_2_M2F_16_net_0 ),
        .GPIO_2_M2F_15                ( ICICLE_MSS_GPIO_2_M2F_15 ),
        .GPIO_2_M2F_14                ( ICICLE_MSS_GPIO_2_M2F_14 ),
        .GPIO_2_M2F_13                ( ICICLE_MSS_GPIO_2_M2F_13 ),
        .GPIO_2_M2F_12                ( ICICLE_MSS_GPIO_2_M2F_12 ),
        .GPIO_2_M2F_11                ( ICICLE_MSS_GPIO_2_M2F_11 ),
        .GPIO_2_M2F_10                ( ICICLE_MSS_GPIO_2_M2F_10 ),
        .GPIO_2_M2F_9                 ( ICICLE_MSS_GPIO_2_M2F_9 ),
        .GPIO_2_M2F_8                 ( ICICLE_MSS_GPIO_2_M2F_8 ),
        .GPIO_2_M2F_7                 ( ICICLE_MSS_GPIO_2_M2F_7 ),
        .GPIO_2_M2F_6                 (  ),
        .GPIO_2_M2F_5                 ( ICICLE_MSS_GPIO_2_M2F_5 ),
        .GPIO_2_M2F_4                 ( ICICLE_MSS_GPIO_2_M2F_4 ),
        .GPIO_2_M2F_3                 ( ICICLE_MSS_GPIO_2_M2F_3 ),
        .GPIO_2_M2F_2                 ( ICICLE_MSS_GPIO_2_M2F_2 ),
        .GPIO_2_M2F_1                 (  ),
        .GPIO_2_M2F_0                 (  ),
        .GPIO_2_OE_M2F_15             ( ICICLE_MSS_GPIO_2_OE_M2F_15 ),
        .GPIO_2_OE_M2F_14             ( ICICLE_MSS_GPIO_2_OE_M2F_14 ),
        .GPIO_2_OE_M2F_13             ( ICICLE_MSS_GPIO_2_OE_M2F_13 ),
        .GPIO_2_OE_M2F_12             ( ICICLE_MSS_GPIO_2_OE_M2F_12 ),
        .GPIO_2_OE_M2F_11             ( ICICLE_MSS_GPIO_2_OE_M2F_11 ),
        .GPIO_2_OE_M2F_10             ( ICICLE_MSS_GPIO_2_OE_M2F_10 ),
        .GPIO_2_OE_M2F_9              ( ICICLE_MSS_GPIO_2_OE_M2F_9 ),
        .GPIO_2_OE_M2F_8              ( ICICLE_MSS_GPIO_2_OE_M2F_8 ),
        .GPIO_2_OE_M2F_7              ( ICICLE_MSS_GPIO_2_OE_M2F_7 ),
        .GPIO_2_OE_M2F_6              (  ),
        .GPIO_2_OE_M2F_5              ( ICICLE_MSS_GPIO_2_OE_M2F_5 ),
        .GPIO_2_OE_M2F_4              ( ICICLE_MSS_GPIO_2_OE_M2F_4 ),
        .GPIO_2_OE_M2F_3              ( ICICLE_MSS_GPIO_2_OE_M2F_3 ),
        .GPIO_2_OE_M2F_2              ( ICICLE_MSS_GPIO_2_OE_M2F_2 ),
        .GPIO_2_OE_M2F_1              (  ),
        .GPIO_2_OE_M2F_0              (  ),
        .PLL_CPU_LOCK_M2F             (  ),
        .PLL_DDR_LOCK_M2F             (  ),
        .PLL_SGMII_LOCK_M2F           (  ),
        .MSS_RESET_N_M2F              ( MSS_RESET_N_M2F_net_0 ),
        .MAC_0_TSU_SOF_TX_M2F         (  ),
        .MAC_0_TSU_SYNC_FRAME_TX_M2F  (  ),
        .MAC_0_TSU_DELAY_REQ_TX_M2F   (  ),
        .MAC_0_TSU_PDELAY_REQ_TX_M2F  (  ),
        .MAC_0_TSU_PDELAY_RESP_TX_M2F (  ),
        .MAC_0_TSU_SOF_RX_M2F         (  ),
        .MAC_0_TSU_SYNC_FRAME_RX_M2F  (  ),
        .MAC_0_TSU_DELAY_REQ_RX_M2F   (  ),
        .MAC_0_TSU_PDELAY_REQ_RX_M2F  (  ),
        .MAC_0_TSU_PDELAY_RESP_RX_M2F (  ),
        .MAC_1_TSU_SOF_TX_M2F         (  ),
        .MAC_1_TSU_SYNC_FRAME_TX_M2F  (  ),
        .MAC_1_TSU_DELAY_REQ_TX_M2F   (  ),
        .MAC_1_TSU_PDELAY_REQ_TX_M2F  (  ),
        .MAC_1_TSU_PDELAY_RESP_TX_M2F (  ),
        .MAC_1_TSU_SOF_RX_M2F         (  ),
        .MAC_1_TSU_SYNC_FRAME_RX_M2F  (  ),
        .MAC_1_TSU_DELAY_REQ_RX_M2F   (  ),
        .MAC_1_TSU_PDELAY_REQ_RX_M2F  (  ),
        .MAC_1_TSU_PDELAY_RESP_RX_M2F (  ),
        .CAN_1_TXBUS                  ( CAN_1_TXBUS_net_0 ),
        .CAN_1_TX_EBL_N               ( CAN_1_TX_EBL_N_net_0 ),
        .MAC_1_MDC                    ( MAC_1_MDC_net_0 ),
        .USB_STP                      ( USB_STP_net_0 ),
        .SPI_1_DO                     ( SPI_1_DO_net_0 ),
        .SD_CLK_EMMC_CLK              ( SD_CLK_EMMC_CLK_net_0 ),
        .SD_POW_EMMC_DATA4            ( SD_POW_EMMC_DATA4_net_0 ),
        .SD_VOLT_SEL_EMMC_DATA5       ( SD_VOLT_SEL_EMMC_DATA5_net_0 ),
        .SD_VOLT_EN_EMMC_DATA6        ( SD_VOLT_EN_EMMC_DATA6_net_0 ),
        .SD_VOLT_CMD_DIR_EMMC_DATA7   ( SD_VOLT_CMD_DIR_EMMC_DATA7_net_0 ),
        .SD_VOLT_DIR_0_EMMC_UNUSED    ( SD_VOLT_DIR_0_EMMC_UNUSED_net_0 ),
        .SD_VOLT_DIR_1_3_EMMC_UNUSED  ( SD_VOLT_DIR_1_3_EMMC_UNUSED_net_0 ),
        .SGMII_TX1_P                  ( SGMII_TX1_P_net_0 ),
        .SGMII_TX1_N                  ( SGMII_TX1_N_net_0 ),
        .SGMII_TX0_P                  ( SGMII_TX0_P_net_0 ),
        .SGMII_TX0_N                  ( SGMII_TX0_N_net_0 ),
        .RESET_N                      ( RESET_N_net_0 ),
        .ODT                          ( ODT_net_0 ),
        .CKE                          ( CKE_net_0 ),
        .CS                           ( CS_net_0 ),
        .CK                           ( CK_net_0 ),
        .CK_N                         ( CK_N_net_0 ),
        .FIC_0_AXI4_M_AWID            ( FIC_0_AXI4_INITIATOR_AWID ),
        .FIC_0_AXI4_M_AWADDR          ( FIC_0_AXI4_INITIATOR_AWADDR ),
        .FIC_0_AXI4_M_AWLEN           ( FIC_0_AXI4_INITIATOR_AWLEN ),
        .FIC_0_AXI4_M_AWSIZE          ( FIC_0_AXI4_INITIATOR_AWSIZE ),
        .FIC_0_AXI4_M_AWBURST         ( FIC_0_AXI4_INITIATOR_AWBURST ),
        .FIC_0_AXI4_M_AWQOS           ( FIC_0_AXI4_INITIATOR_AWQOS ),
        .FIC_0_AXI4_M_AWCACHE         ( FIC_0_AXI4_INITIATOR_AWCACHE ),
        .FIC_0_AXI4_M_AWPROT          ( FIC_0_AXI4_INITIATOR_AWPROT ),
        .FIC_0_AXI4_M_WDATA           ( FIC_0_AXI4_INITIATOR_WDATA ),
        .FIC_0_AXI4_M_WSTRB           ( FIC_0_AXI4_INITIATOR_WSTRB ),
        .FIC_0_AXI4_M_ARID            ( FIC_0_AXI4_INITIATOR_ARID ),
        .FIC_0_AXI4_M_ARADDR          ( FIC_0_AXI4_INITIATOR_ARADDR ),
        .FIC_0_AXI4_M_ARLEN           ( FIC_0_AXI4_INITIATOR_ARLEN ),
        .FIC_0_AXI4_M_ARSIZE          ( FIC_0_AXI4_INITIATOR_ARSIZE ),
        .FIC_0_AXI4_M_ARBURST         ( FIC_0_AXI4_INITIATOR_ARBURST ),
        .FIC_0_AXI4_M_ARQOS           ( FIC_0_AXI4_INITIATOR_ARQOS ),
        .FIC_0_AXI4_M_ARCACHE         ( FIC_0_AXI4_INITIATOR_ARCACHE ),
        .FIC_0_AXI4_M_ARPROT          ( FIC_0_AXI4_INITIATOR_ARPROT ),
        .FIC_0_AXI4_S_BID             ( FIC_0_AXI4_TARGET_BID ),
        .FIC_0_AXI4_S_BRESP           ( FIC_0_AXI4_TARGET_BRESP ),
        .FIC_0_AXI4_S_RID             ( FIC_0_AXI4_TARGET_RID ),
        .FIC_0_AXI4_S_RDATA           ( FIC_0_AXI4_TARGET_RDATA ),
        .FIC_0_AXI4_S_RRESP           ( FIC_0_AXI4_TARGET_RRESP ),
        .FIC_1_AXI4_M_AWID            ( FIC_1_AXI4_INITIATOR_AWID ),
        .FIC_1_AXI4_M_AWADDR          ( FIC_1_AXI4_INITIATOR_AWADDR ),
        .FIC_1_AXI4_M_AWLEN           ( FIC_1_AXI4_INITIATOR_AWLEN ),
        .FIC_1_AXI4_M_AWSIZE          ( FIC_1_AXI4_INITIATOR_AWSIZE ),
        .FIC_1_AXI4_M_AWBURST         ( FIC_1_AXI4_INITIATOR_AWBURST ),
        .FIC_1_AXI4_M_AWQOS           ( FIC_1_AXI4_INITIATOR_AWQOS ),
        .FIC_1_AXI4_M_AWCACHE         ( FIC_1_AXI4_INITIATOR_AWCACHE ),
        .FIC_1_AXI4_M_AWPROT          ( FIC_1_AXI4_INITIATOR_AWPROT ),
        .FIC_1_AXI4_M_WDATA           ( FIC_1_AXI4_INITIATOR_WDATA ),
        .FIC_1_AXI4_M_WSTRB           ( FIC_1_AXI4_INITIATOR_WSTRB ),
        .FIC_1_AXI4_M_ARID            ( FIC_1_AXI4_INITIATOR_ARID ),
        .FIC_1_AXI4_M_ARADDR          ( FIC_1_AXI4_INITIATOR_ARADDR ),
        .FIC_1_AXI4_M_ARLEN           ( FIC_1_AXI4_INITIATOR_ARLEN ),
        .FIC_1_AXI4_M_ARSIZE          ( FIC_1_AXI4_INITIATOR_ARSIZE ),
        .FIC_1_AXI4_M_ARBURST         ( FIC_1_AXI4_INITIATOR_ARBURST ),
        .FIC_1_AXI4_M_ARQOS           ( FIC_1_AXI4_INITIATOR_ARQOS ),
        .FIC_1_AXI4_M_ARCACHE         ( FIC_1_AXI4_INITIATOR_ARCACHE ),
        .FIC_1_AXI4_M_ARPROT          ( FIC_1_AXI4_INITIATOR_ARPROT ),
        .FIC_1_AXI4_S_BID             ( FIC_1_AXI4_TARGET_BID ),
        .FIC_1_AXI4_S_BRESP           ( FIC_1_AXI4_TARGET_BRESP ),
        .FIC_1_AXI4_S_RID             ( FIC_1_AXI4_TARGET_RID ),
        .FIC_1_AXI4_S_RDATA           ( FIC_1_AXI4_TARGET_RDATA ),
        .FIC_1_AXI4_S_RRESP           ( FIC_1_AXI4_TARGET_RRESP ),
        .FIC_2_AXI4_S_BID             ( FIC_2_AXI4_TARGET_BID ),
        .FIC_2_AXI4_S_BRESP           ( FIC_2_AXI4_TARGET_BRESP ),
        .FIC_2_AXI4_S_RID             ( FIC_2_AXI4_TARGET_RID ),
        .FIC_2_AXI4_S_RDATA           ( FIC_2_AXI4_TARGET_RDATA ),
        .FIC_2_AXI4_S_RRESP           ( FIC_2_AXI4_TARGET_RRESP ),
        .FIC_3_APB_M_PADDR            ( FIC_3_APB_INITIATOR_PADDR ),
        .FIC_3_APB_M_PSTRB            (  ),
        .FIC_3_APB_M_PWDATA           ( FIC_3_APB_INITIATOR_PWDATA ),
        .QSPI_DATA_M2F                ( QSPI_DATA_M2F_net_0 ),
        .QSPI_DATA_OE_M2F             ( QSPI_DATA_OE_M2F_net_0 ),
        .MSS_INT_M2F                  (  ),
        .DM                           ( DM_net_0 ),
        .CA                           ( CA_net_0 ),
        // Inouts
        .I2C_1_SCL                    ( I2C_1_SCL ),
        .I2C_1_SDA                    ( I2C_1_SDA ),
        .MAC_1_MDIO                   ( MAC_1_MDIO ),
        .USB_DATA0                    ( USB_DATA0 ),
        .USB_DATA1                    ( USB_DATA1 ),
        .USB_DATA2                    ( USB_DATA2 ),
        .USB_DATA3                    ( USB_DATA3 ),
        .USB_DATA4                    ( USB_DATA4 ),
        .USB_DATA5                    ( USB_DATA5 ),
        .USB_DATA6                    ( USB_DATA6 ),
        .USB_DATA7                    ( USB_DATA7 ),
        .SPI_1_SS0                    ( SPI_1_SS0 ),
        .SPI_1_CLK                    ( SPI_1_CLK ),
        .SD_CMD_EMMC_CMD              ( SD_CMD_EMMC_CMD ),
        .SD_DATA0_EMMC_DATA0          ( SD_DATA0_EMMC_DATA0 ),
        .SD_DATA1_EMMC_DATA1          ( SD_DATA1_EMMC_DATA1 ),
        .SD_DATA2_EMMC_DATA2          ( SD_DATA2_EMMC_DATA2 ),
        .SD_DATA3_EMMC_DATA3          ( SD_DATA3_EMMC_DATA3 ),
        .DQ                           ( DQ ),
        .DQS                          ( DQS ),
        .DQS_N                        ( DQS_N ) 
        );

//--------BIBUF
BIBUF QSPI_CLK_BIBUF(
        // Inputs
        .D   ( ICICLE_MSS_QSPI_CLK_M2F ),
        .E   ( ICICLE_MSS_QSPI_CLK_OE_M2F ),
        // Outputs
        .Y   (  ),
        // Inouts
        .PAD ( QSPI_CLK ) 
        );

//--------BIBUF
BIBUF QSPI_DATA_0_BIBUF(
        // Inputs
        .D   ( ICICLE_MSS_QSPI_DATA_M2F0to0 ),
        .E   ( ICICLE_MSS_QSPI_DATA_OE_M2F0to0 ),
        // Outputs
        .Y   ( QSPI_DATA_0_BIBUF_Y ),
        // Inouts
        .PAD ( QSPI_DATA_0 ) 
        );

//--------BIBUF
BIBUF QSPI_DATA_1_BIBUF(
        // Inputs
        .D   ( ICICLE_MSS_QSPI_DATA_M2F1to1 ),
        .E   ( ICICLE_MSS_QSPI_DATA_OE_M2F1to1 ),
        // Outputs
        .Y   ( QSPI_DATA_1_BIBUF_Y ),
        // Inouts
        .PAD ( QSPI_DATA_1 ) 
        );

//--------BIBUF
BIBUF QSPI_DATA_2_BIBUF(
        // Inputs
        .D   ( ICICLE_MSS_QSPI_DATA_M2F2to2 ),
        .E   ( ICICLE_MSS_QSPI_DATA_OE_M2F2to2 ),
        // Outputs
        .Y   ( QSPI_DATA_2_BIBUF_Y ),
        // Inouts
        .PAD ( QSPI_DATA_2 ) 
        );

//--------BIBUF
BIBUF QSPI_DATA_3_BIBUF(
        // Inputs
        .D   ( ICICLE_MSS_QSPI_DATA_M2F3to3 ),
        .E   ( ICICLE_MSS_QSPI_DATA_OE_M2F3to3 ),
        // Outputs
        .Y   ( QSPI_DATA_3_BIBUF_Y ),
        // Inouts
        .PAD ( QSPI_DATA_3 ) 
        );

//--------BIBUF
BIBUF QSPI_SEL_BIBUF(
        // Inputs
        .D   ( ICICLE_MSS_QSPI_SEL_M2F ),
        .E   ( ICICLE_MSS_QSPI_SEL_OE_M2F ),
        // Outputs
        .Y   (  ),
        // Inouts
        .PAD ( QSPI_SEL ) 
        );


endmodule
