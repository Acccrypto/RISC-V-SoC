///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: tf_ROM.v
// File history:
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// <Description here>
//
// Targeted device: <Family::PolarFireSoC> <Die::MPFS250T_ES> <Package::FCVG484>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

//`timescale <time_units> / <precision>

module tf0_ROM (
    input                       clk,
    input      [5:0]            A,
    output reg [22:0]           Q
);
    
    always@(posedge clk) begin
        case(A)
            6'd0: Q <= 23'd4808194;
            6'd1: Q <= 23'd3765607;
            6'd2: Q <= 23'd3761513;
            6'd3: Q <= 23'd5178923;
            6'd4: Q <= 23'd5496691;
            6'd5: Q <= 23'd5234739;
            6'd6: Q <= 23'd5178987;
            6'd7: Q <= 23'd7778734;
            6'd8: Q <= 23'd3542485;
            6'd9: Q <= 23'd2682288;
            6'd10: Q <= 23'd2129892;
            6'd11: Q <= 23'd3764867;
            6'd12: Q <= 23'd7375178;
            6'd13: Q <= 23'd557458;
            6'd14: Q <= 23'd7159240;
            6'd15: Q <= 23'd5010068;
            6'd16: Q <= 23'd4317364;
            6'd17: Q <= 23'd2663378;
            6'd18: Q <= 23'd6705802;
            6'd19: Q <= 23'd4855975;
            6'd20: Q <= 23'd7946292;
            6'd21: Q <= 23'd676590;
            6'd22: Q <= 23'd7044481;
            6'd23: Q <= 23'd5152541;
            6'd24: Q <= 23'd1714295;
            6'd25: Q <= 23'd2453983;
            6'd26: Q <= 23'd1460718;
            6'd27: Q <= 23'd7737789;
            6'd28: Q <= 23'd4795319;
            6'd29: Q <= 23'd2815639;
            6'd30: Q <= 23'd2283733;
            6'd31: Q <= 23'd3602218;
            6'd32: Q <= 23'd3182878;
            6'd33: Q <= 23'd2740543;
            6'd34: Q <= 23'd4793971;
            6'd35: Q <= 23'd5269599;
            6'd36: Q <= 23'd2101410;
            6'd37: Q <= 23'd3704823;
            6'd38: Q <= 23'd1159875;
            6'd39: Q <= 23'd394148;
            6'd40: Q <= 23'd928749;
            6'd41: Q <= 23'd1095468;
            6'd42: Q <= 23'd4874037;
            6'd43: Q <= 23'd2071829;
            6'd44: Q <= 23'd4361428;
            6'd45: Q <= 23'd3241972;
            6'd46: Q <= 23'd2156050;
            6'd47: Q <= 23'd3415069;
            6'd48: Q <= 23'd1759347;
            6'd49: Q <= 23'd7562881;
            6'd50: Q <= 23'd4805951;
            6'd51: Q <= 23'd3756790;
            6'd52: Q <= 23'd6444618;
            6'd53: Q <= 23'd6663429;
            6'd54: Q <= 23'd4430364;
            6'd55: Q <= 23'd5483103;
            6'd56: Q <= 23'd3192354;
            6'd57: Q <= 23'd556856;
            6'd58: Q <= 23'd3870317;
            6'd59: Q <= 23'd2917338;
            6'd60: Q <= 23'd1853806;
            6'd61: Q <= 23'd3345963;
            6'd62: Q <= 23'd1858416;
        endcase  
    end
    
endmodule
    
module tf1_ROM (
    input                       clk,
    input      [4:0]            A,
    output reg [45:0]           Q
);
    
    always@(posedge clk) begin
        case(A)
            5'd0: Q <= 46'b0101110111000111111000100100110111111010111001;
            5'd1: Q <= 46'b1010111101010010011000001110101100011011101111;
            5'd2: Q <= 46'b0111111110101010100110010011101011001011101010;
            5'd3: Q <= 46'b1010000001111101110000111110111011000101110101;
            5'd4: Q <= 46'b0100110010010001011010000111101111001001010110;
            5'd5: Q <= 46'b0011101100100001010001010001011010011011010100;
            5'd6: Q <= 46'b0101010111001011001101110100100101100010011100;
            5'd7: Q <= 46'b1101110111100011111010101111110111001010001000;
            5'd8: Q <= 46'b0010111010100010000001000001110101110101011001;
            5'd9: Q <= 46'b0010001100001111011101010100101010110010101001;
            5'd10: Q <= 46'b1110111001111101001111000000101001011011011000;
            5'd11: Q <= 46'b0100101100100101110110010011001111111100010010;
            5'd12: Q <= 46'b1000000010011001110100010010101010010110000010;
            5'd13: Q <= 46'b0011110010101001110011010011110001011011000001;
            5'd14: Q <= 46'b0011010011111100111100100000111001011110001111;
            5'd15: Q <= 46'b1001110010010000001011101100011011100001011001;
            5'd16: Q <= 46'b1011000100001001100110000110110100100000100111;
            5'd17: Q <= 46'b1011011011000111101000010111010111100001111010;
            5'd18: Q <= 46'b0110101001000100101111010000000000110001111110;
            5'd19: Q <= 46'b1101100000010011101000110110111101010100110010;
            5'd20: Q <= 46'b1101011110001001101001101001011000111011001011;
            5'd21: Q <= 46'b0101110010100110100110000010010111101001101100;
            5'd22: Q <= 46'b0111011100010000010000011011010010100001011100;
            5'd23: Q <= 46'b0101100101001001111100001100110111110010101010;
            5'd24: Q <= 46'b0010100101100101010000010101011000010100110110;
            5'd25: Q <= 46'b0101000111100011000011010101010111100101011101;
            5'd26: Q <= 46'b1001010111101100111000001000110100101010000110;
            5'd27: Q <= 46'b1110101111010000010011011110001101111001100110;
            5'd28: Q <= 46'b0000101010100101000110011110101101111101011001;
            5'd29: Q <= 46'b0001111011011100001011110110111111001111011010;
            5'd30: Q <= 46'b1000101100110110111111011000101000101100110100;
            5'd31: Q <= 46'b1011101101111101100101100110101001111001111011;
        endcase  
    end

endmodule

module tf2_ROM (
    input                       clk,
    input      [4:0]            A,
    output reg [91:0]           Q
);
    
    always@(posedge clk) begin
        case(A)
            5'd0: Q <= 92'b00000000000011011011001110001001010111110001011010111010010110011110011010011010100011101111;
            5'd1: Q <= 92'b01010001001100000111000110010010110101111111101111110111110001111010101010100100111001111000;
            5'd2: Q <= 92'b00100100000101000100011000000101010100101010000001001101101111111111110000110101111010000111;
            5'd3: Q <= 92'b10000110111111111111000101110011010101101101001001101110000000100111010001110010100010101111;
            5'd4: Q <= 92'b11111110111001101011101000110010001101000011010001111011001101101010110110100110110110000000;
            5'd5: Q <= 92'b11000011010101110011000001100001011101100101101000011011111110011000110001101000001010011000;
            5'd6: Q <= 92'b11001100010100101100000100101111010101011110010101000110111100000011010001100101110110001101;
            5'd7: Q <= 92'b10010011011000011100011000100110110100001101001111100000011011011001110110100110100010110000;
            5'd8: Q <= 92'b10000001001101110101001110010011010011110101010100001011101100010101011001011000010110010001;
            5'd9: Q <= 92'b01001000110111000111001100100011000011100110111111011110001110101100110011110101100001011001;
            5'd10: Q <= 92'b01110010010110110110010010001100001001001000110010010111010110110011110001010100110111110010;
            5'd11: Q <= 92'b01100001100001100011100010100001010100001001000010011001000110010111011111111010111110000000;
            5'd12: Q <= 92'b01011011011111111001011000001000101010000010111111110100000110010110001001100101100001111010;
            5'd13: Q <= 92'b11010110011001101110101000100101011011011101101101011111000011100110010111100000011000011110;
            5'd14: Q <= 92'b11110001110000000001101110001010001100001101110111101101001100000010010010101110010100111100;
            5'd15: Q <= 92'b00111110001110101101000110001100110000101110111110011011000011011100010111101010000001101100;
            5'd16: Q <= 92'b11001110001101011000111010000000011111110001101011011101001001111111111000001101011101110010;
            5'd17: Q <= 92'b00010001111001000000001110110111100000001001000001000000011100110110110101100000001110001110;
            5'd18: Q <= 92'b11010010101011010001000001111001101101001111100100110000000111011110111010101001110111111010;
            5'd19: Q <= 92'b00001111100000000010111110110110111111110101001110100110100001011110111000111110000111100011;
            5'd20: Q <= 92'b10100011001010101110011111101010110110000011010101000011001111011101001011011110110011010100;
            5'd21: Q <= 92'b10110000000000110001100011111101001100111101010001011011100000000100110000100111111000100011;
            5'd22: Q <= 92'b01111001011110100110111010011100110011001100111100111001110010101011100110100100101101011101;
            5'd23: Q <= 92'b00110010110100100100110001111011110010000001100010001110000010100111010011000111011011001000;
            5'd24: Q <= 92'b01111001111010000101111111111110110001100110101101010111101100110110001011100001011001101001;
            5'd25: Q <= 92'b01100110101001011010110000001101000111011000000001000010100100110000011101000001111001111000;
            5'd26: Q <= 92'b01011110110001100010110110111100001010000100010000111110000001111000111101110110110100001011;
            5'd27: Q <= 92'b00011010001111111110000011010001011000001001000000010001000111101010011010001100010101011001;
            5'd28: Q <= 92'b10111101000100010000101010111110101010001100100100011111111000110010110111100110100101000010;
            5'd29: Q <= 92'b10100011110000011101101110010110101101101100110101100101001011110011011110011110000111111110;
            5'd30: Q <= 92'b11110110100000001100100011010111100001110111011000011001110101010110010001100100101011011110;
            5'd31: Q <= 92'b00111001111111000010100111001111110001110011100010000000101110000111011101001011011011010111;
        endcase  
    end

endmodule

