`timescale 1 ns/100 ps
// Version: 


module MSS(
       FIC_0_ACLK,
       FIC_0_AXI4_M_AWREADY,
       FIC_0_AXI4_M_WREADY,
       FIC_0_AXI4_M_BID,
       FIC_0_AXI4_M_BRESP,
       FIC_0_AXI4_M_BVALID,
       FIC_0_AXI4_M_ARREADY,
       FIC_0_AXI4_M_RID,
       FIC_0_AXI4_M_RDATA,
       FIC_0_AXI4_M_RRESP,
       FIC_0_AXI4_M_RLAST,
       FIC_0_AXI4_M_RVALID,
       FIC_0_AXI4_S_AWID,
       FIC_0_AXI4_S_AWADDR,
       FIC_0_AXI4_S_AWLEN,
       FIC_0_AXI4_S_AWSIZE,
       FIC_0_AXI4_S_AWBURST,
       FIC_0_AXI4_S_AWQOS,
       FIC_0_AXI4_S_AWLOCK,
       FIC_0_AXI4_S_AWCACHE,
       FIC_0_AXI4_S_AWPROT,
       FIC_0_AXI4_S_AWVALID,
       FIC_0_AXI4_S_WDATA,
       FIC_0_AXI4_S_WSTRB,
       FIC_0_AXI4_S_WLAST,
       FIC_0_AXI4_S_WVALID,
       FIC_0_AXI4_S_BREADY,
       FIC_0_AXI4_S_ARID,
       FIC_0_AXI4_S_ARADDR,
       FIC_0_AXI4_S_ARLEN,
       FIC_0_AXI4_S_ARSIZE,
       FIC_0_AXI4_S_ARBURST,
       FIC_0_AXI4_S_ARQOS,
       FIC_0_AXI4_S_ARLOCK,
       FIC_0_AXI4_S_ARCACHE,
       FIC_0_AXI4_S_ARPROT,
       FIC_0_AXI4_S_ARVALID,
       FIC_0_AXI4_S_RREADY,
       FIC_1_ACLK,
       FIC_1_AXI4_M_AWREADY,
       FIC_1_AXI4_M_WREADY,
       FIC_1_AXI4_M_BID,
       FIC_1_AXI4_M_BRESP,
       FIC_1_AXI4_M_BVALID,
       FIC_1_AXI4_M_ARREADY,
       FIC_1_AXI4_M_RID,
       FIC_1_AXI4_M_RDATA,
       FIC_1_AXI4_M_RRESP,
       FIC_1_AXI4_M_RLAST,
       FIC_1_AXI4_M_RVALID,
       FIC_1_AXI4_S_AWID,
       FIC_1_AXI4_S_AWADDR,
       FIC_1_AXI4_S_AWLEN,
       FIC_1_AXI4_S_AWSIZE,
       FIC_1_AXI4_S_AWBURST,
       FIC_1_AXI4_S_AWLOCK,
       FIC_1_AXI4_S_AWCACHE,
       FIC_1_AXI4_S_AWQOS,
       FIC_1_AXI4_S_AWPROT,
       FIC_1_AXI4_S_AWVALID,
       FIC_1_AXI4_S_WDATA,
       FIC_1_AXI4_S_WSTRB,
       FIC_1_AXI4_S_WLAST,
       FIC_1_AXI4_S_WVALID,
       FIC_1_AXI4_S_BREADY,
       FIC_1_AXI4_S_ARID,
       FIC_1_AXI4_S_ARADDR,
       FIC_1_AXI4_S_ARLEN,
       FIC_1_AXI4_S_ARSIZE,
       FIC_1_AXI4_S_ARBURST,
       FIC_1_AXI4_S_ARQOS,
       FIC_1_AXI4_S_ARLOCK,
       FIC_1_AXI4_S_ARCACHE,
       FIC_1_AXI4_S_ARPROT,
       FIC_1_AXI4_S_ARVALID,
       FIC_1_AXI4_S_RREADY,
       FIC_2_ACLK,
       SPARE_3_F2M,
       FIC_2_AXI4_S_AWID,
       FIC_2_AXI4_S_AWADDR,
       FIC_2_AXI4_S_AWLEN,
       FIC_2_AXI4_S_AWSIZE,
       FIC_2_AXI4_S_AWBURST,
       FIC_2_AXI4_S_AWLOCK,
       FIC_2_AXI4_S_AWCACHE,
       FIC_2_AXI4_S_AWQOS,
       FIC_2_AXI4_S_AWPROT,
       FIC_2_AXI4_S_AWVALID,
       FIC_2_AXI4_S_WDATA,
       FIC_2_AXI4_S_WSTRB,
       FIC_2_AXI4_S_WLAST,
       FIC_2_AXI4_S_WVALID,
       FIC_2_AXI4_S_BREADY,
       FIC_2_AXI4_S_ARID,
       FIC_2_AXI4_S_ARADDR,
       FIC_2_AXI4_S_ARLEN,
       FIC_2_AXI4_S_ARSIZE,
       FIC_2_AXI4_S_ARBURST,
       FIC_2_AXI4_S_ARLOCK,
       FIC_2_AXI4_S_ARCACHE,
       FIC_2_AXI4_S_ARQOS,
       FIC_2_AXI4_S_ARPROT,
       FIC_2_AXI4_S_ARVALID,
       FIC_2_AXI4_S_RREADY,
       FIC_3_PCLK,
       SPARE_4_F2M,
       FIC_3_APB_M_PRDATA,
       FIC_3_APB_M_PREADY,
       FIC_3_APB_M_PSLVERR,
       MMUART_0_DCD_F2M,
       MMUART_0_RI_F2M,
       MMUART_0_DSR_F2M,
       MMUART_0_CTS_F2M,
       MMUART_0_RXD_F2M,
       MMUART_0_CLK_F2M,
       MMUART_1_DCD_F2M,
       MMUART_1_RI_F2M,
       MMUART_1_DSR_F2M,
       MMUART_1_CTS_F2M,
       MMUART_1_RXD_F2M,
       MMUART_1_CLK_F2M,
       MMUART_2_RXD_F2M,
       MMUART_3_RXD_F2M,
       MMUART_4_RXD_F2M,
       CAN_0_RXBUS_F2M,
       CAN_1_RXBUS_F2M,
       CAN_CLK_F2M,
       QSPI_DATA_F2M,
       SPI_0_SS_F2M,
       SPI_0_DI_F2M,
       SPI_0_CLK_F2M,
       SPI_1_SS_F2M,
       SPI_1_DI_F2M,
       SPI_1_CLK_F2M,
       I2C_0_SCL_F2M,
       I2C_1_SCL_F2M,
       I2C_0_SDA_F2M,
       I2C_1_SDA_F2M,
       I2C_0_BCLK_F2M,
       I2C_0_SMBALERT_NI_F2M,
       I2C_0_SMBSUS_NI_F2M,
       I2C_1_BCLK_F2M,
       I2C_1_SMBALERT_NI_F2M,
       I2C_1_SMBSUS_NI_F2M,
       GPIO_2_F2M,
       MAC_0_MDI_F2M,
       MAC_1_MDI_F2M,
       JTAG_TMS_F2M,
       JTAG_TCK_F2M,
       JTAG_TDI_F2M,
       JTAG_TRSTB_F2M,
       MSS_INT_F2M,
       SPARE_1_F2M,
       SPARE_2_F2M,
       BOOT_FAIL_CLEAR_F2M,
       MSS_RESET_N_F2M,
       GPIO_RESET_N_F2M,
       USOC_TRACE_CLOCK_F2M,
       USOC_TRACE_VALID_F2M,
       USOC_TRACE_DATA_F2M,
       SPARE_5_F2M,
       MAC_0_GMII_MII_RXD_F2M,
       MAC_0_GMII_MII_RX_DV_F2M,
       MAC_0_GMII_MII_RX_ER_F2M,
       MAC_0_GMII_MII_RX_CRS_F2M,
       MAC_0_GMII_MII_RX_COL_F2M,
       MAC_0_GMII_MII_RX_CLK_F2M,
       MAC_0_GMII_MII_TX_CLK_F2M,
       MAC_0_TSU_CLK_F2M,
       MAC_1_GMII_MII_RXD_F2M,
       MAC_1_GMII_MII_RX_DV_F2M,
       MAC_1_GMII_MII_RX_ER_F2M,
       MAC_1_GMII_MII_RX_CRS_F2M,
       MAC_1_GMII_MII_RX_COL_F2M,
       MAC_1_GMII_MII_RX_CLK_F2M,
       MAC_1_GMII_MII_TX_CLK_F2M,
       MAC_1_TSU_CLK_F2M,
       MAC_0_FILTER_MATCH1_F2M,
       MAC_0_FILTER_MATCH2_F2M,
       MAC_0_FILTER_MATCH3_F2M,
       MAC_0_FILTER_MATCH4_F2M,
       MAC_1_FILTER_MATCH1_F2M,
       MAC_1_FILTER_MATCH2_F2M,
       MAC_1_FILTER_MATCH3_F2M,
       MAC_1_FILTER_MATCH4_F2M,
       MAC_0_TSU_GEM_MS_F2M,
       MAC_0_TSU_GEM_INC_CTRL_F2M,
       MAC_1_TSU_GEM_MS_F2M,
       MAC_1_TSU_GEM_INC_CTRL_F2M,
       CRYPTO_HCLK,
       CRYPTO_HRESETN,
       CRYPTO_AHB_M_HREADY,
       CRYPTO_AHB_M_HRESP,
       CRYPTO_AHB_M_HRDATA,
       CRYPTO_AHB_S_HSEL,
       CRYPTO_AHB_S_HADDR,
       CRYPTO_AHB_S_HWDATA,
       CRYPTO_AHB_S_HSIZE,
       CRYPTO_AHB_S_HTRANS,
       CRYPTO_AHB_S_HWRITE,
       CRYPTO_AHB_S_HREADY,
       CRYPTO_STALL_F2M,
       CRYPTO_PURGE_F2M,
       CRYPTO_GO_F2M,
       CRYPTO_REQUEST_F2M,
       CRYPTO_RELEASE_F2M,
       CRYPTO_XENABLE_F2M,
       CRYPTO_XWDATA_F2M,
       CRYPTO_XOUTACK_F2M,
       CRYPTO_MESH_CLEAR_F2M,
       EMMC_SD_CLK_F2M,
       FIC_0_DLL_LOCK_M2F,
       FIC_1_DLL_LOCK_M2F,
       FIC_2_DLL_LOCK_M2F,
       FIC_3_DLL_LOCK_M2F,
       FIC_0_AXI4_M_AWID,
       FIC_0_AXI4_M_AWADDR,
       FIC_0_AXI4_M_AWLEN,
       FIC_0_AXI4_M_AWSIZE,
       FIC_0_AXI4_M_AWBURST,
       FIC_0_AXI4_M_AWLOCK,
       FIC_0_AXI4_M_AWQOS,
       FIC_0_AXI4_M_AWCACHE,
       FIC_0_AXI4_M_AWPROT,
       FIC_0_AXI4_M_AWVALID,
       FIC_0_AXI4_M_WDATA,
       FIC_0_AXI4_M_WSTRB,
       FIC_0_AXI4_M_WLAST,
       FIC_0_AXI4_M_WVALID,
       FIC_0_AXI4_M_BREADY,
       FIC_0_AXI4_M_ARID,
       FIC_0_AXI4_M_ARADDR,
       FIC_0_AXI4_M_ARLEN,
       FIC_0_AXI4_M_ARSIZE,
       FIC_0_AXI4_M_ARBURST,
       FIC_0_AXI4_M_ARLOCK,
       FIC_0_AXI4_M_ARQOS,
       FIC_0_AXI4_M_ARCACHE,
       FIC_0_AXI4_M_ARPROT,
       FIC_0_AXI4_M_ARVALID,
       FIC_0_AXI4_M_RREADY,
       FIC_0_AXI4_S_AWREADY,
       FIC_0_AXI4_S_WREADY,
       FIC_0_AXI4_S_BID,
       FIC_0_AXI4_S_BRESP,
       FIC_0_AXI4_S_BVALID,
       FIC_0_AXI4_S_ARREADY,
       FIC_0_AXI4_S_RID,
       FIC_0_AXI4_S_RDATA,
       FIC_0_AXI4_S_RRESP,
       FIC_0_AXI4_S_RLAST,
       FIC_0_AXI4_S_RVALID,
       FIC_1_AXI4_M_AWID,
       FIC_1_AXI4_M_AWADDR,
       FIC_1_AXI4_M_AWLEN,
       FIC_1_AXI4_M_AWSIZE,
       FIC_1_AXI4_M_AWBURST,
       FIC_1_AXI4_M_AWLOCK,
       FIC_1_AXI4_M_AWQOS,
       FIC_1_AXI4_M_AWCACHE,
       FIC_1_AXI4_M_AWPROT,
       FIC_1_AXI4_M_AWVALID,
       FIC_1_AXI4_M_WDATA,
       FIC_1_AXI4_M_WSTRB,
       FIC_1_AXI4_M_WLAST,
       FIC_1_AXI4_M_WVALID,
       FIC_1_AXI4_M_BREADY,
       FIC_1_AXI4_M_ARID,
       FIC_1_AXI4_M_ARADDR,
       FIC_1_AXI4_M_ARLEN,
       FIC_1_AXI4_M_ARSIZE,
       FIC_1_AXI4_M_ARBURST,
       FIC_1_AXI4_M_ARLOCK,
       FIC_1_AXI4_M_ARQOS,
       FIC_1_AXI4_M_ARCACHE,
       FIC_1_AXI4_M_ARPROT,
       FIC_1_AXI4_M_ARVALID,
       FIC_1_AXI4_M_RREADY,
       FIC_1_AXI4_S_AWREADY,
       FIC_1_AXI4_S_WREADY,
       FIC_1_AXI4_S_BID,
       FIC_1_AXI4_S_BRESP,
       FIC_1_AXI4_S_BVALID,
       FIC_1_AXI4_S_ARREADY,
       FIC_1_AXI4_S_RID,
       FIC_1_AXI4_S_RDATA,
       FIC_1_AXI4_S_RRESP,
       FIC_1_AXI4_S_RLAST,
       FIC_1_AXI4_S_RVALID,
       FIC_2_AXI4_S_AWREADY,
       FIC_2_AXI4_S_WREADY,
       FIC_2_AXI4_S_BID,
       FIC_2_AXI4_S_BRESP,
       FIC_2_AXI4_S_BVALID,
       FIC_2_AXI4_S_ARREADY,
       FIC_2_AXI4_S_RID,
       FIC_2_AXI4_S_RDATA,
       FIC_2_AXI4_S_RRESP,
       FIC_2_AXI4_S_RLAST,
       FIC_2_AXI4_S_RVALID,
       FIC_3_APB_M_PSEL,
       FIC_3_APB_M_PADDR,
       FIC_3_APB_M_PWRITE,
       FIC_3_APB_M_PENABLE,
       FIC_3_APB_M_PSTRB,
       FIC_3_APB_M_PWDATA,
       MMUART_0_DTR_M2F,
       MMUART_0_RTS_M2F,
       MMUART_0_TXD_M2F,
       MMUART_0_TXD_OE_M2F,
       MMUART_1_DTR_M2F,
       MMUART_1_RTS_M2F,
       MMUART_1_TXD_M2F,
       MMUART_1_TXD_OE_M2F,
       MMUART_0_OUT1N_M2F,
       MMUART_0_OUT2N_M2F,
       MMUART_0_TE_M2F,
       MMUART_0_ESWM_M2F,
       MMUART_0_CLK_M2F,
       MMUART_0_CLK_OE_M2F,
       MMUART_1_OUT1N_M2F,
       MMUART_1_OUT2N_M2F,
       MMUART_1_TE_M2F,
       MMUART_1_ESWM_M2F,
       MMUART_1_CLK_M2F,
       MMUART_1_CLK_OE_M2F,
       MMUART_2_TXD_M2F,
       MMUART_3_TXD_M2F,
       MMUART_4_TXD_M2F,
       CAN_0_TX_EBL_M2F,
       CAN_0_TXBUS_M2F,
       CAN_1_TX_EBL_M2F,
       CAN_1_TXBUS_M2F,
       QSPI_SEL_M2F,
       QSPI_SEL_OE_M2F,
       QSPI_CLK_M2F,
       QSPI_CLK_OE_M2F,
       QSPI_DATA_M2F,
       QSPI_DATA_OE_M2F,
       SPI_0_SS1_M2F,
       SPI_0_SS1_OE_M2F,
       SPI_1_SS1_M2F,
       SPI_1_SS1_OE_M2F,
       SPI_0_DO_M2F,
       SPI_0_DO_OE_M2F,
       SPI_0_CLK_M2F,
       SPI_0_CLK_OE_M2F,
       SPI_1_DO_M2F,
       SPI_1_DO_OE_M2F,
       SPI_1_CLK_M2F,
       SPI_1_CLK_OE_M2F,
       I2C_0_SCL_OE_M2F,
       I2C_0_SDA_OE_M2F,
       I2C_1_SCL_OE_M2F,
       I2C_1_SDA_OE_M2F,
       I2C_0_SMBALERT_NO_M2F,
       I2C_0_SMBSUS_NO_M2F,
       I2C_1_SMBALERT_NO_M2F,
       I2C_1_SMBSUS_NO_M2F,
       GPIO_2_M2F,
       GPIO_2_OE_M2F,
       MAC_0_MDO_M2F,
       MAC_0_MDO_OE_M2F,
       MAC_0_MDC_M2F,
       MAC_1_MDO_M2F,
       MAC_1_MDO_OE_M2F,
       MAC_1_MDC_M2F,
       JTAG_TDO_M2F,
       JTAG_TDO_OE_M2F,
       MSS_INT_M2F,
       SPARE_M2F,
       PLL_CPU_LOCK_M2F,
       PLL_DDR_LOCK_M2F,
       PLL_SGMII_LOCK_M2F,
       MSS_STATUS_M2F,
       BOOT_FAIL_ERROR_M2F,
       MSS_RESET_N_M2F,
       SPARE_2_M2F,
       SPARE_3_M2F,
       SPARE_4_M2F,
       SPARE_5_M2F,
       WDOG_0_INTERRUPT_M2F,
       WDOG_1_INTERRUPT_M2F,
       WDOG_2_INTERRUPT_M2F,
       WDOG_3_INTERRUPT_M2F,
       WDOG_4_INTERRUPT_M2F,
       MPU_VIOLATION_FROM_FIC_0_M2F,
       MPU_VIOLATION_FROM_FIC_1_M2F,
       MPU_VIOLATION_FROM_FIC_2_M2F,
       MPU_VIOLATION_FROM_CRYPTO_M2F,
       MPU_VIOLATION_FROM_MAC_0_M2F,
       MPU_VIOLATION_FROM_MAC_1_M2F,
       MPU_VIOLATION_FROM_USB_M2F,
       MPU_VIOLATION_FROM_EMMC_SD_M2F,
       MPU_VIOLATION_FROM_SCB_M2F,
       MPU_VIOLATION_FROM_TRACE_M2F,
       REBOOT_REQUESTED_M2F,
       CPU_IN_RESET_M2F,
       AXI_IN_RESET_M2F,
       SCB_PERIPH_RESET_OCCURRED_M2F,
       SCB_MSS_RESET_OCCURRED_M2F,
       SCB_CPU_RESET_OCCURRED_M2F,
       DEBUGGER_RESET_OCCURRED_M2F,
       FABRIC_RESET_OCCURRED_M2F,
       WDOG_RESET_OCCURRED_M2F,
       GPIO_RESET_OCCURRED_M2F,
       SCB_BUS_RESET_OCCURRED_M2F,
       CPU_SOFT_RESET_OCCURRED_M2F,
       CPU_CLK_DIVIDER_M2F,
       AXI_CLK_DIVIDER_M2F,
       AHB_APB_CLK_DIVIDER_M2F,
       USOC_CONTROL_DATA_M2F,
       MAC_0_GMII_MII_TXD_M2F,
       MAC_0_GMII_MII_TX_EN_M2F,
       MAC_0_GMII_MII_TX_ER_M2F,
       MAC_0_LOCAL_LOOPBACK_M2F,
       MAC_0_LOOPBACK_M2F,
       MAC_0_HALF_DUPLEX_M2F,
       MAC_0_SPEED_MODE_M2F,
       MAC_1_GMII_MII_TXD_M2F,
       MAC_1_GMII_MII_TX_EN_M2F,
       MAC_1_GMII_MII_TX_ER_M2F,
       MAC_1_LOCAL_LOOPBACK_M2F,
       MAC_1_LOOPBACK_M2F,
       MAC_1_HALF_DUPLEX_M2F,
       MAC_1_SPEED_MODE_M2F,
       MAC_0_FILTER_DATA_M2F,
       MAC_0_FILTER_SA_STB_M2F,
       MAC_0_FILTER_DA_STB_M2F,
       MAC_0_FILTER_TYPE_STB_M2F,
       MAC_0_FILTER_VLAN_TAG1_STB_M2F,
       MAC_0_FILTER_VLAN_TAG2_STB_M2F,
       MAC_0_FILTER_IP_SA_STB_M2F,
       MAC_0_FILTER_IP_DA_STB_M2F,
       MAC_0_FILTER_SP_STB_M2F,
       MAC_0_FILTER_DP_STB_M2F,
       MAC_0_FILTER_IPV6_M2F,
       MAC_0_WOL_M2F,
       MAC_1_FILTER_DATA_M2F,
       MAC_1_FILTER_SA_STB_M2F,
       MAC_1_FILTER_DA_STB_M2F,
       MAC_1_FILTER_TYPE_STB_M2F,
       MAC_1_FILTER_VLAN_TAG1_STB_M2F,
       MAC_1_FILTER_VLAN_TAG2_STB_M2F,
       MAC_1_FILTER_IP_SA_STB_M2F,
       MAC_1_FILTER_IP_DA_STB_M2F,
       MAC_1_FILTER_SP_STB_M2F,
       MAC_1_FILTER_DP_STB_M2F,
       MAC_1_FILTER_IPV6_M2F,
       MAC_1_WOL_M2F,
       MAC_0_TSU_SOF_TX_M2F,
       MAC_0_TSU_SYNC_FRAME_TX_M2F,
       MAC_0_TSU_DELAY_REQ_TX_M2F,
       MAC_0_TSU_PDELAY_REQ_TX_M2F,
       MAC_0_TSU_PDELAY_RESP_TX_M2F,
       MAC_0_TSU_SOF_RX_M2F,
       MAC_0_TSU_SYNC_FRAME_RX_M2F,
       MAC_0_TSU_DELAY_REQ_RX_M2F,
       MAC_0_TSU_PDELAY_REQ_RX_M2F,
       MAC_0_TSU_PDELAY_RESP_RX_M2F,
       MAC_0_TSU_TIMER_CNT_M2F,
       MAC_0_TSU_TIMER_CMP_VAL_M2F,
       MAC_1_TSU_SOF_TX_M2F,
       MAC_1_TSU_SYNC_FRAME_TX_M2F,
       MAC_1_TSU_DELAY_REQ_TX_M2F,
       MAC_1_TSU_PDELAY_REQ_TX_M2F,
       MAC_1_TSU_PDELAY_RESP_TX_M2F,
       MAC_1_TSU_SOF_RX_M2F,
       MAC_1_TSU_SYNC_FRAME_RX_M2F,
       MAC_1_TSU_DELAY_REQ_RX_M2F,
       MAC_1_TSU_PDELAY_REQ_RX_M2F,
       MAC_1_TSU_PDELAY_RESP_RX_M2F,
       MAC_1_TSU_TIMER_CNT_M2F,
       MAC_1_TSU_TIMER_CMP_VAL_M2F,
       CRYPTO_DLL_LOCK_M2F,
       CRYPTO_AHB_M_HADDR,
       CRYPTO_AHB_M_HWDATA,
       CRYPTO_AHB_M_HSIZE,
       CRYPTO_AHB_M_HTRANS,
       CRYPTO_AHB_M_HWRITE,
       CRYPTO_AHB_M_HMASTLOCK,
       CRYPTO_AHB_S_HREADYOUT,
       CRYPTO_AHB_S_HRESP,
       CRYPTO_AHB_S_HRDATA,
       CRYPTO_BUSY_M2F,
       CRYPTO_COMPLETE_M2F,
       CRYPTO_ALARM_M2F,
       CRYPTO_BUSERROR_M2F,
       CRYPTO_MSS_REQUEST_M2F,
       CRYPTO_MSS_RELEASE_M2F,
       CRYPTO_OWNER_M2F,
       CRYPTO_MSS_OWNER_M2F,
       CRYPTO_XWADDR_M2F,
       CRYPTO_XINACCEPT_M2F,
       CRYPTO_XRDATA_M2F,
       CRYPTO_XRADDR_M2F,
       CRYPTO_XVALIDOUT_M2F,
       CRYPTO_MESH_ERROR_M2F,
       MSSIO37_IN,
       MSSIO37_OUT,
       MSSIO37_OE,
       MSSIO36_IN,
       MSSIO36_OUT,
       MSSIO36_OE,
       MSSIO35_IN,
       MSSIO35_OUT,
       MSSIO35_OE,
       MSSIO34_IN,
       MSSIO34_OUT,
       MSSIO34_OE,
       MSSIO33_IN,
       MSSIO33_OUT,
       MSSIO33_OE,
       MSSIO32_IN,
       MSSIO32_OUT,
       MSSIO32_OE,
       MSSIO31_IN,
       MSSIO31_OUT,
       MSSIO31_OE,
       MSSIO30_IN,
       MSSIO30_OUT,
       MSSIO30_OE,
       MSSIO29_IN,
       MSSIO29_OUT,
       MSSIO29_OE,
       MSSIO28_IN,
       MSSIO28_OUT,
       MSSIO28_OE,
       MSSIO27_IN,
       MSSIO27_OUT,
       MSSIO27_OE,
       MSSIO26_IN,
       MSSIO26_OUT,
       MSSIO26_OE,
       MSSIO25_IN,
       MSSIO25_OUT,
       MSSIO25_OE,
       MSSIO24_IN,
       MSSIO24_OUT,
       MSSIO24_OE,
       MSSIO23_IN,
       MSSIO23_OUT,
       MSSIO23_OE,
       MSSIO22_IN,
       MSSIO22_OUT,
       MSSIO22_OE,
       MSSIO21_IN,
       MSSIO21_OUT,
       MSSIO21_OE,
       MSSIO20_IN,
       MSSIO20_OUT,
       MSSIO20_OE,
       MSSIO19_IN,
       MSSIO19_OUT,
       MSSIO19_OE,
       MSSIO18_IN,
       MSSIO18_OUT,
       MSSIO18_OE,
       MSSIO17_IN,
       MSSIO17_OUT,
       MSSIO17_OE,
       MSSIO16_IN,
       MSSIO16_OUT,
       MSSIO16_OE,
       MSSIO15_IN,
       MSSIO15_OUT,
       MSSIO15_OE,
       MSSIO14_IN,
       MSSIO14_OUT,
       MSSIO14_OE,
       MSSIO13_IN,
       MSSIO13_OUT,
       MSSIO13_OE,
       MSSIO12_IN,
       MSSIO12_OUT,
       MSSIO12_OE,
       MSSIO11_IN,
       MSSIO11_OUT,
       MSSIO11_OE,
       MSSIO10_IN,
       MSSIO10_OUT,
       MSSIO10_OE,
       MSSIO9_IN,
       MSSIO9_OUT,
       MSSIO9_OE,
       MSSIO8_IN,
       MSSIO8_OUT,
       MSSIO8_OE,
       MSSIO7_IN,
       MSSIO7_OUT,
       MSSIO7_OE,
       MSSIO6_IN,
       MSSIO6_OUT,
       MSSIO6_OE,
       MSSIO5_IN,
       MSSIO5_OUT,
       MSSIO5_OE,
       MSSIO4_IN,
       MSSIO4_OUT,
       MSSIO4_OE,
       MSSIO3_IN,
       MSSIO3_OUT,
       MSSIO3_OE,
       MSSIO2_IN,
       MSSIO2_OUT,
       MSSIO2_OE,
       MSSIO1_IN,
       MSSIO1_OUT,
       MSSIO1_OE,
       MSSIO0_IN,
       MSSIO0_OUT,
       MSSIO0_OE,
       REFCLK,
       SGMII_RX1,
       SGMII_RX0,
       SGMII_TX1,
       SGMII_TX0,
       DDR_DQS4_IN,
       DDR_DQS4_OUT,
       DDR_DQS4_OE,
       DDR_DQS3_IN,
       DDR_DQS3_OUT,
       DDR_DQS3_OE,
       DDR_DQS2_IN,
       DDR_DQS2_OUT,
       DDR_DQS2_OE,
       DDR_DQS1_IN,
       DDR_DQS1_OUT,
       DDR_DQS1_OE,
       DDR_DQS0_IN,
       DDR_DQS0_OUT,
       DDR_DQS0_OE,
       DDR_CK1,
       DDR_CK0,
       DDR3_WE_N,
       DDR_PARITY,
       DDR_RAM_RST_N,
       DDR_ALERT_N,
       DDR_ACT_N,
       DDR_A16,
       DDR_A15,
       DDR_A14,
       DDR_A13,
       DDR_A12,
       DDR_A11,
       DDR_A10,
       DDR_A9,
       DDR_A8,
       DDR_A7,
       DDR_A6,
       DDR_A5,
       DDR_A4,
       DDR_A3,
       DDR_A2,
       DDR_A1,
       DDR_A0,
       DDR_BA1,
       DDR_BA0,
       DDR_BG1,
       DDR_BG0,
       DDR_CKE1,
       DDR_CKE0,
       DDR_CS1,
       DDR_CS0,
       DDR_ODT1,
       DDR_ODT0,
       DDR_DQ35_IN,
       DDR_DQ35_OUT,
       DDR_DQ35_OE,
       DDR_DQ34_IN,
       DDR_DQ34_OUT,
       DDR_DQ34_OE,
       DDR_DQ33_IN,
       DDR_DQ33_OUT,
       DDR_DQ33_OE,
       DDR_DQ32_IN,
       DDR_DQ32_OUT,
       DDR_DQ32_OE,
       DDR_DQ31_IN,
       DDR_DQ31_OUT,
       DDR_DQ31_OE,
       DDR_DQ30_IN,
       DDR_DQ30_OUT,
       DDR_DQ30_OE,
       DDR_DQ29_IN,
       DDR_DQ29_OUT,
       DDR_DQ29_OE,
       DDR_DQ28_IN,
       DDR_DQ28_OUT,
       DDR_DQ28_OE,
       DDR_DQ27_IN,
       DDR_DQ27_OUT,
       DDR_DQ27_OE,
       DDR_DQ26_IN,
       DDR_DQ26_OUT,
       DDR_DQ26_OE,
       DDR_DQ25_IN,
       DDR_DQ25_OUT,
       DDR_DQ25_OE,
       DDR_DQ24_IN,
       DDR_DQ24_OUT,
       DDR_DQ24_OE,
       DDR_DQ23_IN,
       DDR_DQ23_OUT,
       DDR_DQ23_OE,
       DDR_DQ22_IN,
       DDR_DQ22_OUT,
       DDR_DQ22_OE,
       DDR_DQ21_IN,
       DDR_DQ21_OUT,
       DDR_DQ21_OE,
       DDR_DQ20_IN,
       DDR_DQ20_OUT,
       DDR_DQ20_OE,
       DDR_DQ19_IN,
       DDR_DQ19_OUT,
       DDR_DQ19_OE,
       DDR_DQ18_IN,
       DDR_DQ18_OUT,
       DDR_DQ18_OE,
       DDR_DQ17_IN,
       DDR_DQ17_OUT,
       DDR_DQ17_OE,
       DDR_DQ16_IN,
       DDR_DQ16_OUT,
       DDR_DQ16_OE,
       DDR_DQ15_IN,
       DDR_DQ15_OUT,
       DDR_DQ15_OE,
       DDR_DQ14_IN,
       DDR_DQ14_OUT,
       DDR_DQ14_OE,
       DDR_DQ13_IN,
       DDR_DQ13_OUT,
       DDR_DQ13_OE,
       DDR_DQ12_IN,
       DDR_DQ12_OUT,
       DDR_DQ12_OE,
       DDR_DQ11_IN,
       DDR_DQ11_OUT,
       DDR_DQ11_OE,
       DDR_DQ10_IN,
       DDR_DQ10_OUT,
       DDR_DQ10_OE,
       DDR_DQ9_IN,
       DDR_DQ9_OUT,
       DDR_DQ9_OE,
       DDR_DQ8_IN,
       DDR_DQ8_OUT,
       DDR_DQ8_OE,
       DDR_DQ7_IN,
       DDR_DQ7_OUT,
       DDR_DQ7_OE,
       DDR_DQ6_IN,
       DDR_DQ6_OUT,
       DDR_DQ6_OE,
       DDR_DQ5_IN,
       DDR_DQ5_OUT,
       DDR_DQ5_OE,
       DDR_DQ4_IN,
       DDR_DQ4_OUT,
       DDR_DQ4_OE,
       DDR_DQ3_IN,
       DDR_DQ3_OUT,
       DDR_DQ3_OE,
       DDR_DQ2_IN,
       DDR_DQ2_OUT,
       DDR_DQ2_OE,
       DDR_DQ1_IN,
       DDR_DQ1_OUT,
       DDR_DQ1_OE,
       DDR_DQ0_IN,
       DDR_DQ0_OUT,
       DDR_DQ0_OE,
       DDR_DM0_IN,
       DDR_DM0_OUT,
       DDR_DM0_OE,
       DDR_DM1_IN,
       DDR_DM1_OUT,
       DDR_DM1_OE,
       DDR_DM2_IN,
       DDR_DM2_OUT,
       DDR_DM2_OE,
       DDR_DM3_IN,
       DDR_DM3_OUT,
       DDR_DM3_OE,
       DDR_DM4_IN,
       DDR_DM4_OUT,
       DDR_DM4_OE,
       REFCLK_0_PLL_NW,
       REFCLK_1_PLL_NW
    ) ;
/* synthesis syn_black_box

syn_tsu0 = " CRYPTO_AHB_M_HRDATA[0]->CRYPTO_HCLK = 0"
syn_tsu1 = " CRYPTO_AHB_M_HRDATA[10]->CRYPTO_HCLK = 0"
syn_tsu2 = " CRYPTO_AHB_M_HRDATA[11]->CRYPTO_HCLK = 0"
syn_tsu3 = " CRYPTO_AHB_M_HRDATA[12]->CRYPTO_HCLK = 0"
syn_tsu4 = " CRYPTO_AHB_M_HRDATA[13]->CRYPTO_HCLK = 0"
syn_tsu5 = " CRYPTO_AHB_M_HRDATA[14]->CRYPTO_HCLK = 0"
syn_tsu6 = " CRYPTO_AHB_M_HRDATA[15]->CRYPTO_HCLK = 0"
syn_tsu7 = " CRYPTO_AHB_M_HRDATA[16]->CRYPTO_HCLK = 0"
syn_tsu8 = " CRYPTO_AHB_M_HRDATA[17]->CRYPTO_HCLK = 0"
syn_tsu9 = " CRYPTO_AHB_M_HRDATA[18]->CRYPTO_HCLK = 0"
syn_tsu10 = " CRYPTO_AHB_M_HRDATA[19]->CRYPTO_HCLK = 0"
syn_tsu11 = " CRYPTO_AHB_M_HRDATA[1]->CRYPTO_HCLK = 0"
syn_tsu12 = " CRYPTO_AHB_M_HRDATA[20]->CRYPTO_HCLK = 0"
syn_tsu13 = " CRYPTO_AHB_M_HRDATA[21]->CRYPTO_HCLK = 0"
syn_tsu14 = " CRYPTO_AHB_M_HRDATA[22]->CRYPTO_HCLK = 0.028"
syn_tsu15 = " CRYPTO_AHB_M_HRDATA[23]->CRYPTO_HCLK = 0"
syn_tsu16 = " CRYPTO_AHB_M_HRDATA[24]->CRYPTO_HCLK = 0"
syn_tsu17 = " CRYPTO_AHB_M_HRDATA[25]->CRYPTO_HCLK = 0"
syn_tsu18 = " CRYPTO_AHB_M_HRDATA[26]->CRYPTO_HCLK = 0"
syn_tsu19 = " CRYPTO_AHB_M_HRDATA[27]->CRYPTO_HCLK = 0"
syn_tsu20 = " CRYPTO_AHB_M_HRDATA[28]->CRYPTO_HCLK = 0"
syn_tsu21 = " CRYPTO_AHB_M_HRDATA[29]->CRYPTO_HCLK = 0"
syn_tsu22 = " CRYPTO_AHB_M_HRDATA[2]->CRYPTO_HCLK = 0"
syn_tsu23 = " CRYPTO_AHB_M_HRDATA[30]->CRYPTO_HCLK = 0"
syn_tsu24 = " CRYPTO_AHB_M_HRDATA[31]->CRYPTO_HCLK = 0"
syn_tsu25 = " CRYPTO_AHB_M_HRDATA[3]->CRYPTO_HCLK = 0"
syn_tsu26 = " CRYPTO_AHB_M_HRDATA[4]->CRYPTO_HCLK = 0"
syn_tsu27 = " CRYPTO_AHB_M_HRDATA[5]->CRYPTO_HCLK = 0"
syn_tsu28 = " CRYPTO_AHB_M_HRDATA[6]->CRYPTO_HCLK = 0"
syn_tsu29 = " CRYPTO_AHB_M_HRDATA[7]->CRYPTO_HCLK = 0"
syn_tsu30 = " CRYPTO_AHB_M_HRDATA[8]->CRYPTO_HCLK = 0"
syn_tsu31 = " CRYPTO_AHB_M_HRDATA[9]->CRYPTO_HCLK = 0"
syn_tsu32 = " CRYPTO_AHB_M_HREADY->CRYPTO_HCLK = 0"
syn_tsu33 = " CRYPTO_AHB_M_HRESP->CRYPTO_HCLK = 0"
syn_tsu34 = " CRYPTO_AHB_S_HADDR[10]->CRYPTO_HCLK = 0"
syn_tsu35 = " CRYPTO_AHB_S_HADDR[11]->CRYPTO_HCLK = 0"
syn_tsu36 = " CRYPTO_AHB_S_HADDR[12]->CRYPTO_HCLK = 0"
syn_tsu37 = " CRYPTO_AHB_S_HADDR[13]->CRYPTO_HCLK = 0"
syn_tsu38 = " CRYPTO_AHB_S_HADDR[14]->CRYPTO_HCLK = 0"
syn_tsu39 = " CRYPTO_AHB_S_HADDR[15]->CRYPTO_HCLK = 0"
syn_tsu40 = " CRYPTO_AHB_S_HADDR[16]->CRYPTO_HCLK = 0"
syn_tsu41 = " CRYPTO_AHB_S_HADDR[2]->CRYPTO_HCLK = 0"
syn_tsu42 = " CRYPTO_AHB_S_HADDR[3]->CRYPTO_HCLK = 0"
syn_tsu43 = " CRYPTO_AHB_S_HADDR[4]->CRYPTO_HCLK = 0"
syn_tsu44 = " CRYPTO_AHB_S_HADDR[5]->CRYPTO_HCLK = 0"
syn_tsu45 = " CRYPTO_AHB_S_HADDR[6]->CRYPTO_HCLK = 0"
syn_tsu46 = " CRYPTO_AHB_S_HADDR[7]->CRYPTO_HCLK = 0"
syn_tsu47 = " CRYPTO_AHB_S_HADDR[8]->CRYPTO_HCLK = 0"
syn_tsu48 = " CRYPTO_AHB_S_HADDR[9]->CRYPTO_HCLK = 0"
syn_tsu49 = " CRYPTO_AHB_S_HREADY->CRYPTO_HCLK = 0"
syn_tsu50 = " CRYPTO_AHB_S_HSEL->CRYPTO_HCLK = 0"
syn_tsu51 = " CRYPTO_AHB_S_HTRANS[1]->CRYPTO_HCLK = 0"
syn_tsu52 = " CRYPTO_AHB_S_HWDATA[0]->CRYPTO_HCLK = 0"
syn_tsu53 = " CRYPTO_AHB_S_HWDATA[10]->CRYPTO_HCLK = 0"
syn_tsu54 = " CRYPTO_AHB_S_HWDATA[11]->CRYPTO_HCLK = 0"
syn_tsu55 = " CRYPTO_AHB_S_HWDATA[12]->CRYPTO_HCLK = 0"
syn_tsu56 = " CRYPTO_AHB_S_HWDATA[13]->CRYPTO_HCLK = 0"
syn_tsu57 = " CRYPTO_AHB_S_HWDATA[14]->CRYPTO_HCLK = 0"
syn_tsu58 = " CRYPTO_AHB_S_HWDATA[15]->CRYPTO_HCLK = 0"
syn_tsu59 = " CRYPTO_AHB_S_HWDATA[16]->CRYPTO_HCLK = 0"
syn_tsu60 = " CRYPTO_AHB_S_HWDATA[17]->CRYPTO_HCLK = 0"
syn_tsu61 = " CRYPTO_AHB_S_HWDATA[18]->CRYPTO_HCLK = 0"
syn_tsu62 = " CRYPTO_AHB_S_HWDATA[19]->CRYPTO_HCLK = 0"
syn_tsu63 = " CRYPTO_AHB_S_HWDATA[1]->CRYPTO_HCLK = 0"
syn_tsu64 = " CRYPTO_AHB_S_HWDATA[20]->CRYPTO_HCLK = 0"
syn_tsu65 = " CRYPTO_AHB_S_HWDATA[21]->CRYPTO_HCLK = 0"
syn_tsu66 = " CRYPTO_AHB_S_HWDATA[22]->CRYPTO_HCLK = 0"
syn_tsu67 = " CRYPTO_AHB_S_HWDATA[23]->CRYPTO_HCLK = 0"
syn_tsu68 = " CRYPTO_AHB_S_HWDATA[24]->CRYPTO_HCLK = 0"
syn_tsu69 = " CRYPTO_AHB_S_HWDATA[25]->CRYPTO_HCLK = 0"
syn_tsu70 = " CRYPTO_AHB_S_HWDATA[26]->CRYPTO_HCLK = 0"
syn_tsu71 = " CRYPTO_AHB_S_HWDATA[27]->CRYPTO_HCLK = 0"
syn_tsu72 = " CRYPTO_AHB_S_HWDATA[28]->CRYPTO_HCLK = 0"
syn_tsu73 = " CRYPTO_AHB_S_HWDATA[29]->CRYPTO_HCLK = 0"
syn_tsu74 = " CRYPTO_AHB_S_HWDATA[2]->CRYPTO_HCLK = 0"
syn_tsu75 = " CRYPTO_AHB_S_HWDATA[30]->CRYPTO_HCLK = 0"
syn_tsu76 = " CRYPTO_AHB_S_HWDATA[31]->CRYPTO_HCLK = 0"
syn_tsu77 = " CRYPTO_AHB_S_HWDATA[3]->CRYPTO_HCLK = 0"
syn_tsu78 = " CRYPTO_AHB_S_HWDATA[4]->CRYPTO_HCLK = 0"
syn_tsu79 = " CRYPTO_AHB_S_HWDATA[5]->CRYPTO_HCLK = 0"
syn_tsu80 = " CRYPTO_AHB_S_HWDATA[6]->CRYPTO_HCLK = 0"
syn_tsu81 = " CRYPTO_AHB_S_HWDATA[7]->CRYPTO_HCLK = 0"
syn_tsu82 = " CRYPTO_AHB_S_HWDATA[8]->CRYPTO_HCLK = 0"
syn_tsu83 = " CRYPTO_AHB_S_HWDATA[9]->CRYPTO_HCLK = 0"
syn_tsu84 = " CRYPTO_AHB_S_HWRITE->CRYPTO_HCLK = 0"
syn_tsu85 = " CRYPTO_STALL_F2M->CRYPTO_HCLK = 0"
syn_tsu86 = " CRYPTO_XENABLE_F2M->CRYPTO_HCLK = 0"
syn_tsu87 = " CRYPTO_XOUTACK_F2M->CRYPTO_HCLK = 0"
syn_tsu88 = " CRYPTO_XWDATA_F2M[0]->CRYPTO_HCLK = 0"
syn_tsu89 = " CRYPTO_XWDATA_F2M[10]->CRYPTO_HCLK = 0"
syn_tsu90 = " CRYPTO_XWDATA_F2M[11]->CRYPTO_HCLK = 0"
syn_tsu91 = " CRYPTO_XWDATA_F2M[12]->CRYPTO_HCLK = 0"
syn_tsu92 = " CRYPTO_XWDATA_F2M[13]->CRYPTO_HCLK = 0"
syn_tsu93 = " CRYPTO_XWDATA_F2M[14]->CRYPTO_HCLK = 0"
syn_tsu94 = " CRYPTO_XWDATA_F2M[15]->CRYPTO_HCLK = 0"
syn_tsu95 = " CRYPTO_XWDATA_F2M[16]->CRYPTO_HCLK = 0"
syn_tsu96 = " CRYPTO_XWDATA_F2M[17]->CRYPTO_HCLK = 0"
syn_tsu97 = " CRYPTO_XWDATA_F2M[18]->CRYPTO_HCLK = 0"
syn_tsu98 = " CRYPTO_XWDATA_F2M[19]->CRYPTO_HCLK = 0"
syn_tsu99 = " CRYPTO_XWDATA_F2M[1]->CRYPTO_HCLK = 0"
syn_tsu100 = " CRYPTO_XWDATA_F2M[20]->CRYPTO_HCLK = 0"
syn_tsu101 = " CRYPTO_XWDATA_F2M[21]->CRYPTO_HCLK = 0"
syn_tsu102 = " CRYPTO_XWDATA_F2M[22]->CRYPTO_HCLK = 0"
syn_tsu103 = " CRYPTO_XWDATA_F2M[23]->CRYPTO_HCLK = 0"
syn_tsu104 = " CRYPTO_XWDATA_F2M[24]->CRYPTO_HCLK = 0"
syn_tsu105 = " CRYPTO_XWDATA_F2M[25]->CRYPTO_HCLK = 0"
syn_tsu106 = " CRYPTO_XWDATA_F2M[26]->CRYPTO_HCLK = 0"
syn_tsu107 = " CRYPTO_XWDATA_F2M[27]->CRYPTO_HCLK = 0"
syn_tsu108 = " CRYPTO_XWDATA_F2M[28]->CRYPTO_HCLK = 0"
syn_tsu109 = " CRYPTO_XWDATA_F2M[29]->CRYPTO_HCLK = 0"
syn_tsu110 = " CRYPTO_XWDATA_F2M[2]->CRYPTO_HCLK = 0"
syn_tsu111 = " CRYPTO_XWDATA_F2M[30]->CRYPTO_HCLK = 0"
syn_tsu112 = " CRYPTO_XWDATA_F2M[31]->CRYPTO_HCLK = 0"
syn_tsu113 = " CRYPTO_XWDATA_F2M[3]->CRYPTO_HCLK = 0"
syn_tsu114 = " CRYPTO_XWDATA_F2M[4]->CRYPTO_HCLK = 0"
syn_tsu115 = " CRYPTO_XWDATA_F2M[5]->CRYPTO_HCLK = 0"
syn_tsu116 = " CRYPTO_XWDATA_F2M[6]->CRYPTO_HCLK = 0"
syn_tsu117 = " CRYPTO_XWDATA_F2M[7]->CRYPTO_HCLK = 0"
syn_tsu118 = " CRYPTO_XWDATA_F2M[8]->CRYPTO_HCLK = 0"
syn_tsu119 = " CRYPTO_XWDATA_F2M[9]->CRYPTO_HCLK = 0"
syn_tsu120 = " FIC_0_AXI4_M_ARREADY->FIC_0_ACLK = 0.934"
syn_tsu121 = " FIC_0_AXI4_M_AWREADY->FIC_0_ACLK = 0.948"
syn_tsu122 = " FIC_0_AXI4_M_BID[0]->FIC_0_ACLK = 0.706"
syn_tsu123 = " FIC_0_AXI4_M_BID[1]->FIC_0_ACLK = 0.686"
syn_tsu124 = " FIC_0_AXI4_M_BID[2]->FIC_0_ACLK = 0.669"
syn_tsu125 = " FIC_0_AXI4_M_BID[3]->FIC_0_ACLK = 0.664"
syn_tsu126 = " FIC_0_AXI4_M_BID[4]->FIC_0_ACLK = 0.69"
syn_tsu127 = " FIC_0_AXI4_M_BID[5]->FIC_0_ACLK = 0.658"
syn_tsu128 = " FIC_0_AXI4_M_BID[6]->FIC_0_ACLK = 0.702"
syn_tsu129 = " FIC_0_AXI4_M_BID[7]->FIC_0_ACLK = 0.685"
syn_tsu130 = " FIC_0_AXI4_M_BRESP[0]->FIC_0_ACLK = 0.743"
syn_tsu131 = " FIC_0_AXI4_M_BRESP[1]->FIC_0_ACLK = 0.744"
syn_tsu132 = " FIC_0_AXI4_M_BVALID->FIC_0_ACLK = 0.952"
syn_tsu133 = " FIC_0_AXI4_M_RDATA[0]->FIC_0_ACLK = 1.044"
syn_tsu134 = " FIC_0_AXI4_M_RDATA[10]->FIC_0_ACLK = 1.003"
syn_tsu135 = " FIC_0_AXI4_M_RDATA[11]->FIC_0_ACLK = 0.929"
syn_tsu136 = " FIC_0_AXI4_M_RDATA[12]->FIC_0_ACLK = 0.997"
syn_tsu137 = " FIC_0_AXI4_M_RDATA[13]->FIC_0_ACLK = 0.996"
syn_tsu138 = " FIC_0_AXI4_M_RDATA[14]->FIC_0_ACLK = 1.035"
syn_tsu139 = " FIC_0_AXI4_M_RDATA[15]->FIC_0_ACLK = 0.984"
syn_tsu140 = " FIC_0_AXI4_M_RDATA[16]->FIC_0_ACLK = 1.001"
syn_tsu141 = " FIC_0_AXI4_M_RDATA[17]->FIC_0_ACLK = 0.962"
syn_tsu142 = " FIC_0_AXI4_M_RDATA[18]->FIC_0_ACLK = 0.989"
syn_tsu143 = " FIC_0_AXI4_M_RDATA[19]->FIC_0_ACLK = 0.994"
syn_tsu144 = " FIC_0_AXI4_M_RDATA[1]->FIC_0_ACLK = 0.988"
syn_tsu145 = " FIC_0_AXI4_M_RDATA[20]->FIC_0_ACLK = 0.98"
syn_tsu146 = " FIC_0_AXI4_M_RDATA[21]->FIC_0_ACLK = 1.072"
syn_tsu147 = " FIC_0_AXI4_M_RDATA[22]->FIC_0_ACLK = 1.001"
syn_tsu148 = " FIC_0_AXI4_M_RDATA[23]->FIC_0_ACLK = 0.965"
syn_tsu149 = " FIC_0_AXI4_M_RDATA[24]->FIC_0_ACLK = 1.014"
syn_tsu150 = " FIC_0_AXI4_M_RDATA[25]->FIC_0_ACLK = 1.056"
syn_tsu151 = " FIC_0_AXI4_M_RDATA[26]->FIC_0_ACLK = 1.038"
syn_tsu152 = " FIC_0_AXI4_M_RDATA[27]->FIC_0_ACLK = 1.063"
syn_tsu153 = " FIC_0_AXI4_M_RDATA[28]->FIC_0_ACLK = 1.016"
syn_tsu154 = " FIC_0_AXI4_M_RDATA[29]->FIC_0_ACLK = 1.047"
syn_tsu155 = " FIC_0_AXI4_M_RDATA[2]->FIC_0_ACLK = 1.036"
syn_tsu156 = " FIC_0_AXI4_M_RDATA[30]->FIC_0_ACLK = 0.952"
syn_tsu157 = " FIC_0_AXI4_M_RDATA[31]->FIC_0_ACLK = 1.038"
syn_tsu158 = " FIC_0_AXI4_M_RDATA[32]->FIC_0_ACLK = 0.996"
syn_tsu159 = " FIC_0_AXI4_M_RDATA[33]->FIC_0_ACLK = 0.937"
syn_tsu160 = " FIC_0_AXI4_M_RDATA[34]->FIC_0_ACLK = 0.99"
syn_tsu161 = " FIC_0_AXI4_M_RDATA[35]->FIC_0_ACLK = 0.998"
syn_tsu162 = " FIC_0_AXI4_M_RDATA[36]->FIC_0_ACLK = 1.033"
syn_tsu163 = " FIC_0_AXI4_M_RDATA[37]->FIC_0_ACLK = 1.059"
syn_tsu164 = " FIC_0_AXI4_M_RDATA[38]->FIC_0_ACLK = 1.032"
syn_tsu165 = " FIC_0_AXI4_M_RDATA[39]->FIC_0_ACLK = 0.97"
syn_tsu166 = " FIC_0_AXI4_M_RDATA[3]->FIC_0_ACLK = 1.003"
syn_tsu167 = " FIC_0_AXI4_M_RDATA[40]->FIC_0_ACLK = 0.971"
syn_tsu168 = " FIC_0_AXI4_M_RDATA[41]->FIC_0_ACLK = 1.048"
syn_tsu169 = " FIC_0_AXI4_M_RDATA[42]->FIC_0_ACLK = 1.033"
syn_tsu170 = " FIC_0_AXI4_M_RDATA[43]->FIC_0_ACLK = 0.926"
syn_tsu171 = " FIC_0_AXI4_M_RDATA[44]->FIC_0_ACLK = 1.027"
syn_tsu172 = " FIC_0_AXI4_M_RDATA[45]->FIC_0_ACLK = 0.994"
syn_tsu173 = " FIC_0_AXI4_M_RDATA[46]->FIC_0_ACLK = 1.052"
syn_tsu174 = " FIC_0_AXI4_M_RDATA[47]->FIC_0_ACLK = 1.038"
syn_tsu175 = " FIC_0_AXI4_M_RDATA[48]->FIC_0_ACLK = 0.997"
syn_tsu176 = " FIC_0_AXI4_M_RDATA[49]->FIC_0_ACLK = 1.019"
syn_tsu177 = " FIC_0_AXI4_M_RDATA[4]->FIC_0_ACLK = 0.997"
syn_tsu178 = " FIC_0_AXI4_M_RDATA[50]->FIC_0_ACLK = 1.029"
syn_tsu179 = " FIC_0_AXI4_M_RDATA[51]->FIC_0_ACLK = 1.038"
syn_tsu180 = " FIC_0_AXI4_M_RDATA[52]->FIC_0_ACLK = 0.981"
syn_tsu181 = " FIC_0_AXI4_M_RDATA[53]->FIC_0_ACLK = 0.985"
syn_tsu182 = " FIC_0_AXI4_M_RDATA[54]->FIC_0_ACLK = 0.886"
syn_tsu183 = " FIC_0_AXI4_M_RDATA[55]->FIC_0_ACLK = 1.047"
syn_tsu184 = " FIC_0_AXI4_M_RDATA[56]->FIC_0_ACLK = 0.957"
syn_tsu185 = " FIC_0_AXI4_M_RDATA[57]->FIC_0_ACLK = 0.96"
syn_tsu186 = " FIC_0_AXI4_M_RDATA[58]->FIC_0_ACLK = 1.029"
syn_tsu187 = " FIC_0_AXI4_M_RDATA[59]->FIC_0_ACLK = 1.007"
syn_tsu188 = " FIC_0_AXI4_M_RDATA[5]->FIC_0_ACLK = 1.022"
syn_tsu189 = " FIC_0_AXI4_M_RDATA[60]->FIC_0_ACLK = 1.008"
syn_tsu190 = " FIC_0_AXI4_M_RDATA[61]->FIC_0_ACLK = 0.958"
syn_tsu191 = " FIC_0_AXI4_M_RDATA[62]->FIC_0_ACLK = 0.916"
syn_tsu192 = " FIC_0_AXI4_M_RDATA[63]->FIC_0_ACLK = 1.027"
syn_tsu193 = " FIC_0_AXI4_M_RDATA[6]->FIC_0_ACLK = 1.058"
syn_tsu194 = " FIC_0_AXI4_M_RDATA[7]->FIC_0_ACLK = 1.09"
syn_tsu195 = " FIC_0_AXI4_M_RDATA[8]->FIC_0_ACLK = 1"
syn_tsu196 = " FIC_0_AXI4_M_RDATA[9]->FIC_0_ACLK = 1"
syn_tsu197 = " FIC_0_AXI4_M_RID[0]->FIC_0_ACLK = 0.997"
syn_tsu198 = " FIC_0_AXI4_M_RID[1]->FIC_0_ACLK = 1.04"
syn_tsu199 = " FIC_0_AXI4_M_RID[2]->FIC_0_ACLK = 1.054"
syn_tsu200 = " FIC_0_AXI4_M_RID[3]->FIC_0_ACLK = 0.996"
syn_tsu201 = " FIC_0_AXI4_M_RID[4]->FIC_0_ACLK = 1.054"
syn_tsu202 = " FIC_0_AXI4_M_RID[5]->FIC_0_ACLK = 0.957"
syn_tsu203 = " FIC_0_AXI4_M_RID[6]->FIC_0_ACLK = 1.019"
syn_tsu204 = " FIC_0_AXI4_M_RID[7]->FIC_0_ACLK = 1.009"
syn_tsu205 = " FIC_0_AXI4_M_RLAST->FIC_0_ACLK = 1.013"
syn_tsu206 = " FIC_0_AXI4_M_RRESP[0]->FIC_0_ACLK = 1.028"
syn_tsu207 = " FIC_0_AXI4_M_RRESP[1]->FIC_0_ACLK = 0.99"
syn_tsu208 = " FIC_0_AXI4_M_RVALID->FIC_0_ACLK = 1.056"
syn_tsu209 = " FIC_0_AXI4_M_WREADY->FIC_0_ACLK = 1.015"
syn_tsu210 = " FIC_0_AXI4_S_ARADDR[0]->FIC_0_ACLK = 0.855"
syn_tsu211 = " FIC_0_AXI4_S_ARADDR[10]->FIC_0_ACLK = 0.757"
syn_tsu212 = " FIC_0_AXI4_S_ARADDR[11]->FIC_0_ACLK = 0.783"
syn_tsu213 = " FIC_0_AXI4_S_ARADDR[12]->FIC_0_ACLK = 0.775"
syn_tsu214 = " FIC_0_AXI4_S_ARADDR[13]->FIC_0_ACLK = 0.776"
syn_tsu215 = " FIC_0_AXI4_S_ARADDR[14]->FIC_0_ACLK = 0.805"
syn_tsu216 = " FIC_0_AXI4_S_ARADDR[15]->FIC_0_ACLK = 0.815"
syn_tsu217 = " FIC_0_AXI4_S_ARADDR[16]->FIC_0_ACLK = 0.796"
syn_tsu218 = " FIC_0_AXI4_S_ARADDR[17]->FIC_0_ACLK = 0.752"
syn_tsu219 = " FIC_0_AXI4_S_ARADDR[18]->FIC_0_ACLK = 0.774"
syn_tsu220 = " FIC_0_AXI4_S_ARADDR[19]->FIC_0_ACLK = 0.728"
syn_tsu221 = " FIC_0_AXI4_S_ARADDR[1]->FIC_0_ACLK = 0.849"
syn_tsu222 = " FIC_0_AXI4_S_ARADDR[20]->FIC_0_ACLK = 0.709"
syn_tsu223 = " FIC_0_AXI4_S_ARADDR[21]->FIC_0_ACLK = 0.75"
syn_tsu224 = " FIC_0_AXI4_S_ARADDR[22]->FIC_0_ACLK = 0.734"
syn_tsu225 = " FIC_0_AXI4_S_ARADDR[23]->FIC_0_ACLK = 0.748"
syn_tsu226 = " FIC_0_AXI4_S_ARADDR[24]->FIC_0_ACLK = 0.735"
syn_tsu227 = " FIC_0_AXI4_S_ARADDR[25]->FIC_0_ACLK = 0.734"
syn_tsu228 = " FIC_0_AXI4_S_ARADDR[26]->FIC_0_ACLK = 0.746"
syn_tsu229 = " FIC_0_AXI4_S_ARADDR[27]->FIC_0_ACLK = 0.755"
syn_tsu230 = " FIC_0_AXI4_S_ARADDR[28]->FIC_0_ACLK = 0.712"
syn_tsu231 = " FIC_0_AXI4_S_ARADDR[29]->FIC_0_ACLK = 0.724"
syn_tsu232 = " FIC_0_AXI4_S_ARADDR[2]->FIC_0_ACLK = 0.851"
syn_tsu233 = " FIC_0_AXI4_S_ARADDR[30]->FIC_0_ACLK = 0.751"
syn_tsu234 = " FIC_0_AXI4_S_ARADDR[31]->FIC_0_ACLK = 0.748"
syn_tsu235 = " FIC_0_AXI4_S_ARADDR[32]->FIC_0_ACLK = 0.76"
syn_tsu236 = " FIC_0_AXI4_S_ARADDR[33]->FIC_0_ACLK = 0.791"
syn_tsu237 = " FIC_0_AXI4_S_ARADDR[34]->FIC_0_ACLK = 0.8"
syn_tsu238 = " FIC_0_AXI4_S_ARADDR[35]->FIC_0_ACLK = 0.778"
syn_tsu239 = " FIC_0_AXI4_S_ARADDR[36]->FIC_0_ACLK = 0.788"
syn_tsu240 = " FIC_0_AXI4_S_ARADDR[37]->FIC_0_ACLK = 0.795"
syn_tsu241 = " FIC_0_AXI4_S_ARADDR[3]->FIC_0_ACLK = 0.776"
syn_tsu242 = " FIC_0_AXI4_S_ARADDR[4]->FIC_0_ACLK = 0.771"
syn_tsu243 = " FIC_0_AXI4_S_ARADDR[5]->FIC_0_ACLK = 0.802"
syn_tsu244 = " FIC_0_AXI4_S_ARADDR[6]->FIC_0_ACLK = 0.797"
syn_tsu245 = " FIC_0_AXI4_S_ARADDR[7]->FIC_0_ACLK = 0.766"
syn_tsu246 = " FIC_0_AXI4_S_ARADDR[8]->FIC_0_ACLK = 0.805"
syn_tsu247 = " FIC_0_AXI4_S_ARADDR[9]->FIC_0_ACLK = 0.791"
syn_tsu248 = " FIC_0_AXI4_S_ARBURST[0]->FIC_0_ACLK = 0.915"
syn_tsu249 = " FIC_0_AXI4_S_ARBURST[1]->FIC_0_ACLK = 0.888"
syn_tsu250 = " FIC_0_AXI4_S_ARCACHE[0]->FIC_0_ACLK = 0.858"
syn_tsu251 = " FIC_0_AXI4_S_ARCACHE[1]->FIC_0_ACLK = 0.874"
syn_tsu252 = " FIC_0_AXI4_S_ARCACHE[2]->FIC_0_ACLK = 0.913"
syn_tsu253 = " FIC_0_AXI4_S_ARCACHE[3]->FIC_0_ACLK = 0.883"
syn_tsu254 = " FIC_0_AXI4_S_ARID[0]->FIC_0_ACLK = 0.756"
syn_tsu255 = " FIC_0_AXI4_S_ARID[1]->FIC_0_ACLK = 0.769"
syn_tsu256 = " FIC_0_AXI4_S_ARID[2]->FIC_0_ACLK = 0.756"
syn_tsu257 = " FIC_0_AXI4_S_ARID[3]->FIC_0_ACLK = 0.756"
syn_tsu258 = " FIC_0_AXI4_S_ARLEN[0]->FIC_0_ACLK = 0.817"
syn_tsu259 = " FIC_0_AXI4_S_ARLEN[1]->FIC_0_ACLK = 0.749"
syn_tsu260 = " FIC_0_AXI4_S_ARLEN[2]->FIC_0_ACLK = 0.731"
syn_tsu261 = " FIC_0_AXI4_S_ARLEN[3]->FIC_0_ACLK = 0.736"
syn_tsu262 = " FIC_0_AXI4_S_ARLEN[4]->FIC_0_ACLK = 0.89"
syn_tsu263 = " FIC_0_AXI4_S_ARLEN[5]->FIC_0_ACLK = 0.818"
syn_tsu264 = " FIC_0_AXI4_S_ARLEN[6]->FIC_0_ACLK = 0.786"
syn_tsu265 = " FIC_0_AXI4_S_ARLEN[7]->FIC_0_ACLK = 0.794"
syn_tsu266 = " FIC_0_AXI4_S_ARLOCK->FIC_0_ACLK = 0.685"
syn_tsu267 = " FIC_0_AXI4_S_ARPROT[0]->FIC_0_ACLK = 0.702"
syn_tsu268 = " FIC_0_AXI4_S_ARPROT[1]->FIC_0_ACLK = 0.781"
syn_tsu269 = " FIC_0_AXI4_S_ARPROT[2]->FIC_0_ACLK = 0.78"
syn_tsu270 = " FIC_0_AXI4_S_ARQOS[0]->FIC_0_ACLK = 0.739"
syn_tsu271 = " FIC_0_AXI4_S_ARQOS[1]->FIC_0_ACLK = 0.783"
syn_tsu272 = " FIC_0_AXI4_S_ARQOS[2]->FIC_0_ACLK = 0.78"
syn_tsu273 = " FIC_0_AXI4_S_ARQOS[3]->FIC_0_ACLK = 0.802"
syn_tsu274 = " FIC_0_AXI4_S_ARSIZE[0]->FIC_0_ACLK = 0.704"
syn_tsu275 = " FIC_0_AXI4_S_ARSIZE[1]->FIC_0_ACLK = 0.712"
syn_tsu276 = " FIC_0_AXI4_S_ARSIZE[2]->FIC_0_ACLK = 0.779"
syn_tsu277 = " FIC_0_AXI4_S_ARVALID->FIC_0_ACLK = 1.029"
syn_tsu278 = " FIC_0_AXI4_S_AWADDR[0]->FIC_0_ACLK = 0.726"
syn_tsu279 = " FIC_0_AXI4_S_AWADDR[10]->FIC_0_ACLK = 0.77"
syn_tsu280 = " FIC_0_AXI4_S_AWADDR[11]->FIC_0_ACLK = 0.774"
syn_tsu281 = " FIC_0_AXI4_S_AWADDR[12]->FIC_0_ACLK = 0.782"
syn_tsu282 = " FIC_0_AXI4_S_AWADDR[13]->FIC_0_ACLK = 0.73"
syn_tsu283 = " FIC_0_AXI4_S_AWADDR[14]->FIC_0_ACLK = 0.818"
syn_tsu284 = " FIC_0_AXI4_S_AWADDR[15]->FIC_0_ACLK = 0.748"
syn_tsu285 = " FIC_0_AXI4_S_AWADDR[16]->FIC_0_ACLK = 0.829"
syn_tsu286 = " FIC_0_AXI4_S_AWADDR[17]->FIC_0_ACLK = 0.709"
syn_tsu287 = " FIC_0_AXI4_S_AWADDR[18]->FIC_0_ACLK = 0.802"
syn_tsu288 = " FIC_0_AXI4_S_AWADDR[19]->FIC_0_ACLK = 0.81"
syn_tsu289 = " FIC_0_AXI4_S_AWADDR[1]->FIC_0_ACLK = 0.728"
syn_tsu290 = " FIC_0_AXI4_S_AWADDR[20]->FIC_0_ACLK = 0.726"
syn_tsu291 = " FIC_0_AXI4_S_AWADDR[21]->FIC_0_ACLK = 0.737"
syn_tsu292 = " FIC_0_AXI4_S_AWADDR[22]->FIC_0_ACLK = 0.697"
syn_tsu293 = " FIC_0_AXI4_S_AWADDR[23]->FIC_0_ACLK = 0.689"
syn_tsu294 = " FIC_0_AXI4_S_AWADDR[24]->FIC_0_ACLK = 0.672"
syn_tsu295 = " FIC_0_AXI4_S_AWADDR[25]->FIC_0_ACLK = 0.689"
syn_tsu296 = " FIC_0_AXI4_S_AWADDR[26]->FIC_0_ACLK = 0.679"
syn_tsu297 = " FIC_0_AXI4_S_AWADDR[27]->FIC_0_ACLK = 0.687"
syn_tsu298 = " FIC_0_AXI4_S_AWADDR[28]->FIC_0_ACLK = 0.694"
syn_tsu299 = " FIC_0_AXI4_S_AWADDR[29]->FIC_0_ACLK = 0.685"
syn_tsu300 = " FIC_0_AXI4_S_AWADDR[2]->FIC_0_ACLK = 0.717"
syn_tsu301 = " FIC_0_AXI4_S_AWADDR[30]->FIC_0_ACLK = 0.689"
syn_tsu302 = " FIC_0_AXI4_S_AWADDR[31]->FIC_0_ACLK = 0.691"
syn_tsu303 = " FIC_0_AXI4_S_AWADDR[32]->FIC_0_ACLK = 0.661"
syn_tsu304 = " FIC_0_AXI4_S_AWADDR[33]->FIC_0_ACLK = 0.73"
syn_tsu305 = " FIC_0_AXI4_S_AWADDR[34]->FIC_0_ACLK = 0.758"
syn_tsu306 = " FIC_0_AXI4_S_AWADDR[35]->FIC_0_ACLK = 0.749"
syn_tsu307 = " FIC_0_AXI4_S_AWADDR[36]->FIC_0_ACLK = 0.749"
syn_tsu308 = " FIC_0_AXI4_S_AWADDR[37]->FIC_0_ACLK = 0.765"
syn_tsu309 = " FIC_0_AXI4_S_AWADDR[3]->FIC_0_ACLK = 0.738"
syn_tsu310 = " FIC_0_AXI4_S_AWADDR[4]->FIC_0_ACLK = 0.733"
syn_tsu311 = " FIC_0_AXI4_S_AWADDR[5]->FIC_0_ACLK = 0.73"
syn_tsu312 = " FIC_0_AXI4_S_AWADDR[6]->FIC_0_ACLK = 0.759"
syn_tsu313 = " FIC_0_AXI4_S_AWADDR[7]->FIC_0_ACLK = 0.733"
syn_tsu314 = " FIC_0_AXI4_S_AWADDR[8]->FIC_0_ACLK = 0.758"
syn_tsu315 = " FIC_0_AXI4_S_AWADDR[9]->FIC_0_ACLK = 0.766"
syn_tsu316 = " FIC_0_AXI4_S_AWBURST[0]->FIC_0_ACLK = 0.747"
syn_tsu317 = " FIC_0_AXI4_S_AWBURST[1]->FIC_0_ACLK = 0.743"
syn_tsu318 = " FIC_0_AXI4_S_AWCACHE[0]->FIC_0_ACLK = 0.745"
syn_tsu319 = " FIC_0_AXI4_S_AWCACHE[1]->FIC_0_ACLK = 0.722"
syn_tsu320 = " FIC_0_AXI4_S_AWCACHE[2]->FIC_0_ACLK = 0.779"
syn_tsu321 = " FIC_0_AXI4_S_AWCACHE[3]->FIC_0_ACLK = 0.791"
syn_tsu322 = " FIC_0_AXI4_S_AWID[0]->FIC_0_ACLK = 0.727"
syn_tsu323 = " FIC_0_AXI4_S_AWID[1]->FIC_0_ACLK = 0.706"
syn_tsu324 = " FIC_0_AXI4_S_AWID[2]->FIC_0_ACLK = 0.727"
syn_tsu325 = " FIC_0_AXI4_S_AWID[3]->FIC_0_ACLK = 0.726"
syn_tsu326 = " FIC_0_AXI4_S_AWLEN[0]->FIC_0_ACLK = 0.72"
syn_tsu327 = " FIC_0_AXI4_S_AWLEN[1]->FIC_0_ACLK = 0.701"
syn_tsu328 = " FIC_0_AXI4_S_AWLEN[2]->FIC_0_ACLK = 0.687"
syn_tsu329 = " FIC_0_AXI4_S_AWLEN[3]->FIC_0_ACLK = 0.672"
syn_tsu330 = " FIC_0_AXI4_S_AWLEN[4]->FIC_0_ACLK = 0.674"
syn_tsu331 = " FIC_0_AXI4_S_AWLEN[5]->FIC_0_ACLK = 0.71"
syn_tsu332 = " FIC_0_AXI4_S_AWLEN[6]->FIC_0_ACLK = 0.662"
syn_tsu333 = " FIC_0_AXI4_S_AWLEN[7]->FIC_0_ACLK = 0.673"
syn_tsu334 = " FIC_0_AXI4_S_AWLOCK->FIC_0_ACLK = 0.683"
syn_tsu335 = " FIC_0_AXI4_S_AWPROT[0]->FIC_0_ACLK = 0.689"
syn_tsu336 = " FIC_0_AXI4_S_AWPROT[1]->FIC_0_ACLK = 0.685"
syn_tsu337 = " FIC_0_AXI4_S_AWPROT[2]->FIC_0_ACLK = 0.72"
syn_tsu338 = " FIC_0_AXI4_S_AWQOS[0]->FIC_0_ACLK = 0.745"
syn_tsu339 = " FIC_0_AXI4_S_AWQOS[1]->FIC_0_ACLK = 0.707"
syn_tsu340 = " FIC_0_AXI4_S_AWQOS[2]->FIC_0_ACLK = 0.704"
syn_tsu341 = " FIC_0_AXI4_S_AWQOS[3]->FIC_0_ACLK = 0.686"
syn_tsu342 = " FIC_0_AXI4_S_AWSIZE[0]->FIC_0_ACLK = 0.663"
syn_tsu343 = " FIC_0_AXI4_S_AWSIZE[1]->FIC_0_ACLK = 0.651"
syn_tsu344 = " FIC_0_AXI4_S_AWSIZE[2]->FIC_0_ACLK = 0.666"
syn_tsu345 = " FIC_0_AXI4_S_AWVALID->FIC_0_ACLK = 0.966"
syn_tsu346 = " FIC_0_AXI4_S_BREADY->FIC_0_ACLK = 1.042"
syn_tsu347 = " FIC_0_AXI4_S_RREADY->FIC_0_ACLK = 1.047"
syn_tsu348 = " FIC_0_AXI4_S_WDATA[0]->FIC_0_ACLK = 0.943"
syn_tsu349 = " FIC_0_AXI4_S_WDATA[10]->FIC_0_ACLK = 0.883"
syn_tsu350 = " FIC_0_AXI4_S_WDATA[11]->FIC_0_ACLK = 0.858"
syn_tsu351 = " FIC_0_AXI4_S_WDATA[12]->FIC_0_ACLK = 0.863"
syn_tsu352 = " FIC_0_AXI4_S_WDATA[13]->FIC_0_ACLK = 0.861"
syn_tsu353 = " FIC_0_AXI4_S_WDATA[14]->FIC_0_ACLK = 0.855"
syn_tsu354 = " FIC_0_AXI4_S_WDATA[15]->FIC_0_ACLK = 0.948"
syn_tsu355 = " FIC_0_AXI4_S_WDATA[16]->FIC_0_ACLK = 0.97"
syn_tsu356 = " FIC_0_AXI4_S_WDATA[17]->FIC_0_ACLK = 0.847"
syn_tsu357 = " FIC_0_AXI4_S_WDATA[18]->FIC_0_ACLK = 0.898"
syn_tsu358 = " FIC_0_AXI4_S_WDATA[19]->FIC_0_ACLK = 0.897"
syn_tsu359 = " FIC_0_AXI4_S_WDATA[1]->FIC_0_ACLK = 0.946"
syn_tsu360 = " FIC_0_AXI4_S_WDATA[20]->FIC_0_ACLK = 0.912"
syn_tsu361 = " FIC_0_AXI4_S_WDATA[21]->FIC_0_ACLK = 0.851"
syn_tsu362 = " FIC_0_AXI4_S_WDATA[22]->FIC_0_ACLK = 0.945"
syn_tsu363 = " FIC_0_AXI4_S_WDATA[23]->FIC_0_ACLK = 0.877"
syn_tsu364 = " FIC_0_AXI4_S_WDATA[24]->FIC_0_ACLK = 0.948"
syn_tsu365 = " FIC_0_AXI4_S_WDATA[25]->FIC_0_ACLK = 0.914"
syn_tsu366 = " FIC_0_AXI4_S_WDATA[26]->FIC_0_ACLK = 0.938"
syn_tsu367 = " FIC_0_AXI4_S_WDATA[27]->FIC_0_ACLK = 0.944"
syn_tsu368 = " FIC_0_AXI4_S_WDATA[28]->FIC_0_ACLK = 0.856"
syn_tsu369 = " FIC_0_AXI4_S_WDATA[29]->FIC_0_ACLK = 0.91"
syn_tsu370 = " FIC_0_AXI4_S_WDATA[2]->FIC_0_ACLK = 0.943"
syn_tsu371 = " FIC_0_AXI4_S_WDATA[30]->FIC_0_ACLK = 0.891"
syn_tsu372 = " FIC_0_AXI4_S_WDATA[31]->FIC_0_ACLK = 0.897"
syn_tsu373 = " FIC_0_AXI4_S_WDATA[32]->FIC_0_ACLK = 0.915"
syn_tsu374 = " FIC_0_AXI4_S_WDATA[33]->FIC_0_ACLK = 0.926"
syn_tsu375 = " FIC_0_AXI4_S_WDATA[34]->FIC_0_ACLK = 0.953"
syn_tsu376 = " FIC_0_AXI4_S_WDATA[35]->FIC_0_ACLK = 0.959"
syn_tsu377 = " FIC_0_AXI4_S_WDATA[36]->FIC_0_ACLK = 0.955"
syn_tsu378 = " FIC_0_AXI4_S_WDATA[37]->FIC_0_ACLK = 0.945"
syn_tsu379 = " FIC_0_AXI4_S_WDATA[38]->FIC_0_ACLK = 0.955"
syn_tsu380 = " FIC_0_AXI4_S_WDATA[39]->FIC_0_ACLK = 0.93"
syn_tsu381 = " FIC_0_AXI4_S_WDATA[3]->FIC_0_ACLK = 1.06"
syn_tsu382 = " FIC_0_AXI4_S_WDATA[40]->FIC_0_ACLK = 0.934"
syn_tsu383 = " FIC_0_AXI4_S_WDATA[41]->FIC_0_ACLK = 0.947"
syn_tsu384 = " FIC_0_AXI4_S_WDATA[42]->FIC_0_ACLK = 0.971"
syn_tsu385 = " FIC_0_AXI4_S_WDATA[43]->FIC_0_ACLK = 0.903"
syn_tsu386 = " FIC_0_AXI4_S_WDATA[44]->FIC_0_ACLK = 1.004"
syn_tsu387 = " FIC_0_AXI4_S_WDATA[45]->FIC_0_ACLK = 0.94"
syn_tsu388 = " FIC_0_AXI4_S_WDATA[46]->FIC_0_ACLK = 0.931"
syn_tsu389 = " FIC_0_AXI4_S_WDATA[47]->FIC_0_ACLK = 0.977"
syn_tsu390 = " FIC_0_AXI4_S_WDATA[48]->FIC_0_ACLK = 0.957"
syn_tsu391 = " FIC_0_AXI4_S_WDATA[49]->FIC_0_ACLK = 0.953"
syn_tsu392 = " FIC_0_AXI4_S_WDATA[4]->FIC_0_ACLK = 1.014"
syn_tsu393 = " FIC_0_AXI4_S_WDATA[50]->FIC_0_ACLK = 0.896"
syn_tsu394 = " FIC_0_AXI4_S_WDATA[51]->FIC_0_ACLK = 0.947"
syn_tsu395 = " FIC_0_AXI4_S_WDATA[52]->FIC_0_ACLK = 0.934"
syn_tsu396 = " FIC_0_AXI4_S_WDATA[53]->FIC_0_ACLK = 0.976"
syn_tsu397 = " FIC_0_AXI4_S_WDATA[54]->FIC_0_ACLK = 0.895"
syn_tsu398 = " FIC_0_AXI4_S_WDATA[55]->FIC_0_ACLK = 0.886"
syn_tsu399 = " FIC_0_AXI4_S_WDATA[56]->FIC_0_ACLK = 0.927"
syn_tsu400 = " FIC_0_AXI4_S_WDATA[57]->FIC_0_ACLK = 0.916"
syn_tsu401 = " FIC_0_AXI4_S_WDATA[58]->FIC_0_ACLK = 0.9"
syn_tsu402 = " FIC_0_AXI4_S_WDATA[59]->FIC_0_ACLK = 0.849"
syn_tsu403 = " FIC_0_AXI4_S_WDATA[5]->FIC_0_ACLK = 0.876"
syn_tsu404 = " FIC_0_AXI4_S_WDATA[60]->FIC_0_ACLK = 0.885"
syn_tsu405 = " FIC_0_AXI4_S_WDATA[61]->FIC_0_ACLK = 0.837"
syn_tsu406 = " FIC_0_AXI4_S_WDATA[62]->FIC_0_ACLK = 0.777"
syn_tsu407 = " FIC_0_AXI4_S_WDATA[63]->FIC_0_ACLK = 0.93"
syn_tsu408 = " FIC_0_AXI4_S_WDATA[6]->FIC_0_ACLK = 0.97"
syn_tsu409 = " FIC_0_AXI4_S_WDATA[7]->FIC_0_ACLK = 0.879"
syn_tsu410 = " FIC_0_AXI4_S_WDATA[8]->FIC_0_ACLK = 0.917"
syn_tsu411 = " FIC_0_AXI4_S_WDATA[9]->FIC_0_ACLK = 0.893"
syn_tsu412 = " FIC_0_AXI4_S_WLAST->FIC_0_ACLK = 1.028"
syn_tsu413 = " FIC_0_AXI4_S_WSTRB[0]->FIC_0_ACLK = 0.967"
syn_tsu414 = " FIC_0_AXI4_S_WSTRB[1]->FIC_0_ACLK = 1.046"
syn_tsu415 = " FIC_0_AXI4_S_WSTRB[2]->FIC_0_ACLK = 1.026"
syn_tsu416 = " FIC_0_AXI4_S_WSTRB[3]->FIC_0_ACLK = 1.008"
syn_tsu417 = " FIC_0_AXI4_S_WSTRB[4]->FIC_0_ACLK = 1.008"
syn_tsu418 = " FIC_0_AXI4_S_WSTRB[5]->FIC_0_ACLK = 0.958"
syn_tsu419 = " FIC_0_AXI4_S_WSTRB[6]->FIC_0_ACLK = 1.047"
syn_tsu420 = " FIC_0_AXI4_S_WSTRB[7]->FIC_0_ACLK = 1.026"
syn_tsu421 = " FIC_0_AXI4_S_WVALID->FIC_0_ACLK = 1.011"
syn_tsu422 = " FIC_1_AXI4_M_ARREADY->FIC_1_ACLK = 1.055"
syn_tsu423 = " FIC_1_AXI4_M_AWREADY->FIC_1_ACLK = 1.046"
syn_tsu424 = " FIC_1_AXI4_M_BID[0]->FIC_1_ACLK = 0.845"
syn_tsu425 = " FIC_1_AXI4_M_BID[1]->FIC_1_ACLK = 0.839"
syn_tsu426 = " FIC_1_AXI4_M_BID[2]->FIC_1_ACLK = 0.916"
syn_tsu427 = " FIC_1_AXI4_M_BID[3]->FIC_1_ACLK = 0.832"
syn_tsu428 = " FIC_1_AXI4_M_BID[4]->FIC_1_ACLK = 0.87"
syn_tsu429 = " FIC_1_AXI4_M_BID[5]->FIC_1_ACLK = 0.859"
syn_tsu430 = " FIC_1_AXI4_M_BID[6]->FIC_1_ACLK = 0.831"
syn_tsu431 = " FIC_1_AXI4_M_BID[7]->FIC_1_ACLK = 0.857"
syn_tsu432 = " FIC_1_AXI4_M_BRESP[0]->FIC_1_ACLK = 0.867"
syn_tsu433 = " FIC_1_AXI4_M_BRESP[1]->FIC_1_ACLK = 0.873"
syn_tsu434 = " FIC_1_AXI4_M_BVALID->FIC_1_ACLK = 1.013"
syn_tsu435 = " FIC_1_AXI4_M_RDATA[0]->FIC_1_ACLK = 0.962"
syn_tsu436 = " FIC_1_AXI4_M_RDATA[10]->FIC_1_ACLK = 0.942"
syn_tsu437 = " FIC_1_AXI4_M_RDATA[11]->FIC_1_ACLK = 0.988"
syn_tsu438 = " FIC_1_AXI4_M_RDATA[12]->FIC_1_ACLK = 1.056"
syn_tsu439 = " FIC_1_AXI4_M_RDATA[13]->FIC_1_ACLK = 1.038"
syn_tsu440 = " FIC_1_AXI4_M_RDATA[14]->FIC_1_ACLK = 1.056"
syn_tsu441 = " FIC_1_AXI4_M_RDATA[15]->FIC_1_ACLK = 0.89"
syn_tsu442 = " FIC_1_AXI4_M_RDATA[16]->FIC_1_ACLK = 1.034"
syn_tsu443 = " FIC_1_AXI4_M_RDATA[17]->FIC_1_ACLK = 0.947"
syn_tsu444 = " FIC_1_AXI4_M_RDATA[18]->FIC_1_ACLK = 0.946"
syn_tsu445 = " FIC_1_AXI4_M_RDATA[19]->FIC_1_ACLK = 0.99"
syn_tsu446 = " FIC_1_AXI4_M_RDATA[1]->FIC_1_ACLK = 0.958"
syn_tsu447 = " FIC_1_AXI4_M_RDATA[20]->FIC_1_ACLK = 1.047"
syn_tsu448 = " FIC_1_AXI4_M_RDATA[21]->FIC_1_ACLK = 0.975"
syn_tsu449 = " FIC_1_AXI4_M_RDATA[22]->FIC_1_ACLK = 0.943"
syn_tsu450 = " FIC_1_AXI4_M_RDATA[23]->FIC_1_ACLK = 0.981"
syn_tsu451 = " FIC_1_AXI4_M_RDATA[24]->FIC_1_ACLK = 1.049"
syn_tsu452 = " FIC_1_AXI4_M_RDATA[25]->FIC_1_ACLK = 0.859"
syn_tsu453 = " FIC_1_AXI4_M_RDATA[26]->FIC_1_ACLK = 0.944"
syn_tsu454 = " FIC_1_AXI4_M_RDATA[27]->FIC_1_ACLK = 0.966"
syn_tsu455 = " FIC_1_AXI4_M_RDATA[28]->FIC_1_ACLK = 0.868"
syn_tsu456 = " FIC_1_AXI4_M_RDATA[29]->FIC_1_ACLK = 0.977"
syn_tsu457 = " FIC_1_AXI4_M_RDATA[2]->FIC_1_ACLK = 1.023"
syn_tsu458 = " FIC_1_AXI4_M_RDATA[30]->FIC_1_ACLK = 0.897"
syn_tsu459 = " FIC_1_AXI4_M_RDATA[31]->FIC_1_ACLK = 0.994"
syn_tsu460 = " FIC_1_AXI4_M_RDATA[32]->FIC_1_ACLK = 0.947"
syn_tsu461 = " FIC_1_AXI4_M_RDATA[33]->FIC_1_ACLK = 0.87"
syn_tsu462 = " FIC_1_AXI4_M_RDATA[34]->FIC_1_ACLK = 0.849"
syn_tsu463 = " FIC_1_AXI4_M_RDATA[35]->FIC_1_ACLK = 0.826"
syn_tsu464 = " FIC_1_AXI4_M_RDATA[36]->FIC_1_ACLK = 0.842"
syn_tsu465 = " FIC_1_AXI4_M_RDATA[37]->FIC_1_ACLK = 0.863"
syn_tsu466 = " FIC_1_AXI4_M_RDATA[38]->FIC_1_ACLK = 0.831"
syn_tsu467 = " FIC_1_AXI4_M_RDATA[39]->FIC_1_ACLK = 0.848"
syn_tsu468 = " FIC_1_AXI4_M_RDATA[3]->FIC_1_ACLK = 1.023"
syn_tsu469 = " FIC_1_AXI4_M_RDATA[40]->FIC_1_ACLK = 0.896"
syn_tsu470 = " FIC_1_AXI4_M_RDATA[41]->FIC_1_ACLK = 0.805"
syn_tsu471 = " FIC_1_AXI4_M_RDATA[42]->FIC_1_ACLK = 0.833"
syn_tsu472 = " FIC_1_AXI4_M_RDATA[43]->FIC_1_ACLK = 0.892"
syn_tsu473 = " FIC_1_AXI4_M_RDATA[44]->FIC_1_ACLK = 0.802"
syn_tsu474 = " FIC_1_AXI4_M_RDATA[45]->FIC_1_ACLK = 0.809"
syn_tsu475 = " FIC_1_AXI4_M_RDATA[46]->FIC_1_ACLK = 0.828"
syn_tsu476 = " FIC_1_AXI4_M_RDATA[47]->FIC_1_ACLK = 0.829"
syn_tsu477 = " FIC_1_AXI4_M_RDATA[48]->FIC_1_ACLK = 0.816"
syn_tsu478 = " FIC_1_AXI4_M_RDATA[49]->FIC_1_ACLK = 0.842"
syn_tsu479 = " FIC_1_AXI4_M_RDATA[4]->FIC_1_ACLK = 0.973"
syn_tsu480 = " FIC_1_AXI4_M_RDATA[50]->FIC_1_ACLK = 0.837"
syn_tsu481 = " FIC_1_AXI4_M_RDATA[51]->FIC_1_ACLK = 0.846"
syn_tsu482 = " FIC_1_AXI4_M_RDATA[52]->FIC_1_ACLK = 0.874"
syn_tsu483 = " FIC_1_AXI4_M_RDATA[53]->FIC_1_ACLK = 0.874"
syn_tsu484 = " FIC_1_AXI4_M_RDATA[54]->FIC_1_ACLK = 0.836"
syn_tsu485 = " FIC_1_AXI4_M_RDATA[55]->FIC_1_ACLK = 0.897"
syn_tsu486 = " FIC_1_AXI4_M_RDATA[56]->FIC_1_ACLK = 0.855"
syn_tsu487 = " FIC_1_AXI4_M_RDATA[57]->FIC_1_ACLK = 0.883"
syn_tsu488 = " FIC_1_AXI4_M_RDATA[58]->FIC_1_ACLK = 0.892"
syn_tsu489 = " FIC_1_AXI4_M_RDATA[59]->FIC_1_ACLK = 0.844"
syn_tsu490 = " FIC_1_AXI4_M_RDATA[5]->FIC_1_ACLK = 0.995"
syn_tsu491 = " FIC_1_AXI4_M_RDATA[60]->FIC_1_ACLK = 0.841"
syn_tsu492 = " FIC_1_AXI4_M_RDATA[61]->FIC_1_ACLK = 0.873"
syn_tsu493 = " FIC_1_AXI4_M_RDATA[62]->FIC_1_ACLK = 0.871"
syn_tsu494 = " FIC_1_AXI4_M_RDATA[63]->FIC_1_ACLK = 0.818"
syn_tsu495 = " FIC_1_AXI4_M_RDATA[6]->FIC_1_ACLK = 0.948"
syn_tsu496 = " FIC_1_AXI4_M_RDATA[7]->FIC_1_ACLK = 0.999"
syn_tsu497 = " FIC_1_AXI4_M_RDATA[8]->FIC_1_ACLK = 1.053"
syn_tsu498 = " FIC_1_AXI4_M_RDATA[9]->FIC_1_ACLK = 1.029"
syn_tsu499 = " FIC_1_AXI4_M_RID[0]->FIC_1_ACLK = 0.977"
syn_tsu500 = " FIC_1_AXI4_M_RID[1]->FIC_1_ACLK = 1.033"
syn_tsu501 = " FIC_1_AXI4_M_RID[2]->FIC_1_ACLK = 1.054"
syn_tsu502 = " FIC_1_AXI4_M_RID[3]->FIC_1_ACLK = 0.955"
syn_tsu503 = " FIC_1_AXI4_M_RID[4]->FIC_1_ACLK = 1.041"
syn_tsu504 = " FIC_1_AXI4_M_RID[5]->FIC_1_ACLK = 0.987"
syn_tsu505 = " FIC_1_AXI4_M_RID[6]->FIC_1_ACLK = 1.016"
syn_tsu506 = " FIC_1_AXI4_M_RID[7]->FIC_1_ACLK = 1.029"
syn_tsu507 = " FIC_1_AXI4_M_RLAST->FIC_1_ACLK = 0.95"
syn_tsu508 = " FIC_1_AXI4_M_RRESP[0]->FIC_1_ACLK = 0.964"
syn_tsu509 = " FIC_1_AXI4_M_RRESP[1]->FIC_1_ACLK = 0.962"
syn_tsu510 = " FIC_1_AXI4_M_RVALID->FIC_1_ACLK = 1.046"
syn_tsu511 = " FIC_1_AXI4_M_WREADY->FIC_1_ACLK = 1.068"
syn_tsu512 = " FIC_1_AXI4_S_ARADDR[0]->FIC_1_ACLK = 0.735"
syn_tsu513 = " FIC_1_AXI4_S_ARADDR[10]->FIC_1_ACLK = 0.792"
syn_tsu514 = " FIC_1_AXI4_S_ARADDR[11]->FIC_1_ACLK = 0.863"
syn_tsu515 = " FIC_1_AXI4_S_ARADDR[12]->FIC_1_ACLK = 0.834"
syn_tsu516 = " FIC_1_AXI4_S_ARADDR[13]->FIC_1_ACLK = 0.792"
syn_tsu517 = " FIC_1_AXI4_S_ARADDR[14]->FIC_1_ACLK = 0.828"
syn_tsu518 = " FIC_1_AXI4_S_ARADDR[15]->FIC_1_ACLK = 0.807"
syn_tsu519 = " FIC_1_AXI4_S_ARADDR[16]->FIC_1_ACLK = 0.801"
syn_tsu520 = " FIC_1_AXI4_S_ARADDR[17]->FIC_1_ACLK = 0.802"
syn_tsu521 = " FIC_1_AXI4_S_ARADDR[18]->FIC_1_ACLK = 0.741"
syn_tsu522 = " FIC_1_AXI4_S_ARADDR[19]->FIC_1_ACLK = 0.819"
syn_tsu523 = " FIC_1_AXI4_S_ARADDR[1]->FIC_1_ACLK = 0.802"
syn_tsu524 = " FIC_1_AXI4_S_ARADDR[20]->FIC_1_ACLK = 0.797"
syn_tsu525 = " FIC_1_AXI4_S_ARADDR[21]->FIC_1_ACLK = 0.81"
syn_tsu526 = " FIC_1_AXI4_S_ARADDR[22]->FIC_1_ACLK = 0.802"
syn_tsu527 = " FIC_1_AXI4_S_ARADDR[23]->FIC_1_ACLK = 0.809"
syn_tsu528 = " FIC_1_AXI4_S_ARADDR[24]->FIC_1_ACLK = 0.817"
syn_tsu529 = " FIC_1_AXI4_S_ARADDR[25]->FIC_1_ACLK = 0.746"
syn_tsu530 = " FIC_1_AXI4_S_ARADDR[26]->FIC_1_ACLK = 0.809"
syn_tsu531 = " FIC_1_AXI4_S_ARADDR[27]->FIC_1_ACLK = 0.775"
syn_tsu532 = " FIC_1_AXI4_S_ARADDR[28]->FIC_1_ACLK = 0.795"
syn_tsu533 = " FIC_1_AXI4_S_ARADDR[29]->FIC_1_ACLK = 0.805"
syn_tsu534 = " FIC_1_AXI4_S_ARADDR[2]->FIC_1_ACLK = 0.72"
syn_tsu535 = " FIC_1_AXI4_S_ARADDR[30]->FIC_1_ACLK = 0.791"
syn_tsu536 = " FIC_1_AXI4_S_ARADDR[31]->FIC_1_ACLK = 0.729"
syn_tsu537 = " FIC_1_AXI4_S_ARADDR[32]->FIC_1_ACLK = 0.744"
syn_tsu538 = " FIC_1_AXI4_S_ARADDR[33]->FIC_1_ACLK = 0.824"
syn_tsu539 = " FIC_1_AXI4_S_ARADDR[34]->FIC_1_ACLK = 0.809"
syn_tsu540 = " FIC_1_AXI4_S_ARADDR[35]->FIC_1_ACLK = 0.821"
syn_tsu541 = " FIC_1_AXI4_S_ARADDR[36]->FIC_1_ACLK = 0.832"
syn_tsu542 = " FIC_1_AXI4_S_ARADDR[37]->FIC_1_ACLK = 0.833"
syn_tsu543 = " FIC_1_AXI4_S_ARADDR[3]->FIC_1_ACLK = 0.809"
syn_tsu544 = " FIC_1_AXI4_S_ARADDR[4]->FIC_1_ACLK = 0.79"
syn_tsu545 = " FIC_1_AXI4_S_ARADDR[5]->FIC_1_ACLK = 0.792"
syn_tsu546 = " FIC_1_AXI4_S_ARADDR[6]->FIC_1_ACLK = 0.778"
syn_tsu547 = " FIC_1_AXI4_S_ARADDR[7]->FIC_1_ACLK = 0.865"
syn_tsu548 = " FIC_1_AXI4_S_ARADDR[8]->FIC_1_ACLK = 0.886"
syn_tsu549 = " FIC_1_AXI4_S_ARADDR[9]->FIC_1_ACLK = 0.793"
syn_tsu550 = " FIC_1_AXI4_S_ARBURST[0]->FIC_1_ACLK = 0.781"
syn_tsu551 = " FIC_1_AXI4_S_ARBURST[1]->FIC_1_ACLK = 0.753"
syn_tsu552 = " FIC_1_AXI4_S_ARCACHE[0]->FIC_1_ACLK = 0.832"
syn_tsu553 = " FIC_1_AXI4_S_ARCACHE[1]->FIC_1_ACLK = 0.769"
syn_tsu554 = " FIC_1_AXI4_S_ARCACHE[2]->FIC_1_ACLK = 0.735"
syn_tsu555 = " FIC_1_AXI4_S_ARCACHE[3]->FIC_1_ACLK = 0.825"
syn_tsu556 = " FIC_1_AXI4_S_ARID[0]->FIC_1_ACLK = 0.756"
syn_tsu557 = " FIC_1_AXI4_S_ARID[1]->FIC_1_ACLK = 0.8"
syn_tsu558 = " FIC_1_AXI4_S_ARID[2]->FIC_1_ACLK = 0.747"
syn_tsu559 = " FIC_1_AXI4_S_ARID[3]->FIC_1_ACLK = 0.766"
syn_tsu560 = " FIC_1_AXI4_S_ARLEN[0]->FIC_1_ACLK = 0.756"
syn_tsu561 = " FIC_1_AXI4_S_ARLEN[1]->FIC_1_ACLK = 0.799"
syn_tsu562 = " FIC_1_AXI4_S_ARLEN[2]->FIC_1_ACLK = 0.806"
syn_tsu563 = " FIC_1_AXI4_S_ARLEN[3]->FIC_1_ACLK = 0.776"
syn_tsu564 = " FIC_1_AXI4_S_ARLEN[4]->FIC_1_ACLK = 0.821"
syn_tsu565 = " FIC_1_AXI4_S_ARLEN[5]->FIC_1_ACLK = 0.756"
syn_tsu566 = " FIC_1_AXI4_S_ARLEN[6]->FIC_1_ACLK = 0.877"
syn_tsu567 = " FIC_1_AXI4_S_ARLEN[7]->FIC_1_ACLK = 0.742"
syn_tsu568 = " FIC_1_AXI4_S_ARLOCK->FIC_1_ACLK = 0.788"
syn_tsu569 = " FIC_1_AXI4_S_ARPROT[0]->FIC_1_ACLK = 0.856"
syn_tsu570 = " FIC_1_AXI4_S_ARPROT[1]->FIC_1_ACLK = 0.734"
syn_tsu571 = " FIC_1_AXI4_S_ARPROT[2]->FIC_1_ACLK = 0.72"
syn_tsu572 = " FIC_1_AXI4_S_ARQOS[0]->FIC_1_ACLK = 0.771"
syn_tsu573 = " FIC_1_AXI4_S_ARQOS[1]->FIC_1_ACLK = 0.748"
syn_tsu574 = " FIC_1_AXI4_S_ARQOS[2]->FIC_1_ACLK = 0.736"
syn_tsu575 = " FIC_1_AXI4_S_ARQOS[3]->FIC_1_ACLK = 0.782"
syn_tsu576 = " FIC_1_AXI4_S_ARSIZE[0]->FIC_1_ACLK = 0.769"
syn_tsu577 = " FIC_1_AXI4_S_ARSIZE[1]->FIC_1_ACLK = 0.791"
syn_tsu578 = " FIC_1_AXI4_S_ARSIZE[2]->FIC_1_ACLK = 0.765"
syn_tsu579 = " FIC_1_AXI4_S_ARVALID->FIC_1_ACLK = 1.053"
syn_tsu580 = " FIC_1_AXI4_S_AWADDR[0]->FIC_1_ACLK = 0.76"
syn_tsu581 = " FIC_1_AXI4_S_AWADDR[10]->FIC_1_ACLK = 0.806"
syn_tsu582 = " FIC_1_AXI4_S_AWADDR[11]->FIC_1_ACLK = 0.752"
syn_tsu583 = " FIC_1_AXI4_S_AWADDR[12]->FIC_1_ACLK = 0.838"
syn_tsu584 = " FIC_1_AXI4_S_AWADDR[13]->FIC_1_ACLK = 0.819"
syn_tsu585 = " FIC_1_AXI4_S_AWADDR[14]->FIC_1_ACLK = 0.77"
syn_tsu586 = " FIC_1_AXI4_S_AWADDR[15]->FIC_1_ACLK = 0.828"
syn_tsu587 = " FIC_1_AXI4_S_AWADDR[16]->FIC_1_ACLK = 0.728"
syn_tsu588 = " FIC_1_AXI4_S_AWADDR[17]->FIC_1_ACLK = 0.821"
syn_tsu589 = " FIC_1_AXI4_S_AWADDR[18]->FIC_1_ACLK = 0.719"
syn_tsu590 = " FIC_1_AXI4_S_AWADDR[19]->FIC_1_ACLK = 0.792"
syn_tsu591 = " FIC_1_AXI4_S_AWADDR[1]->FIC_1_ACLK = 0.75"
syn_tsu592 = " FIC_1_AXI4_S_AWADDR[20]->FIC_1_ACLK = 0.738"
syn_tsu593 = " FIC_1_AXI4_S_AWADDR[21]->FIC_1_ACLK = 0.774"
syn_tsu594 = " FIC_1_AXI4_S_AWADDR[22]->FIC_1_ACLK = 0.787"
syn_tsu595 = " FIC_1_AXI4_S_AWADDR[23]->FIC_1_ACLK = 0.733"
syn_tsu596 = " FIC_1_AXI4_S_AWADDR[24]->FIC_1_ACLK = 0.769"
syn_tsu597 = " FIC_1_AXI4_S_AWADDR[25]->FIC_1_ACLK = 0.809"
syn_tsu598 = " FIC_1_AXI4_S_AWADDR[26]->FIC_1_ACLK = 0.761"
syn_tsu599 = " FIC_1_AXI4_S_AWADDR[27]->FIC_1_ACLK = 0.734"
syn_tsu600 = " FIC_1_AXI4_S_AWADDR[28]->FIC_1_ACLK = 0.763"
syn_tsu601 = " FIC_1_AXI4_S_AWADDR[29]->FIC_1_ACLK = 0.728"
syn_tsu602 = " FIC_1_AXI4_S_AWADDR[2]->FIC_1_ACLK = 0.742"
syn_tsu603 = " FIC_1_AXI4_S_AWADDR[30]->FIC_1_ACLK = 0.735"
syn_tsu604 = " FIC_1_AXI4_S_AWADDR[31]->FIC_1_ACLK = 0.777"
syn_tsu605 = " FIC_1_AXI4_S_AWADDR[32]->FIC_1_ACLK = 0.856"
syn_tsu606 = " FIC_1_AXI4_S_AWADDR[33]->FIC_1_ACLK = 0.818"
syn_tsu607 = " FIC_1_AXI4_S_AWADDR[34]->FIC_1_ACLK = 0.859"
syn_tsu608 = " FIC_1_AXI4_S_AWADDR[35]->FIC_1_ACLK = 0.826"
syn_tsu609 = " FIC_1_AXI4_S_AWADDR[36]->FIC_1_ACLK = 0.782"
syn_tsu610 = " FIC_1_AXI4_S_AWADDR[37]->FIC_1_ACLK = 0.876"
syn_tsu611 = " FIC_1_AXI4_S_AWADDR[3]->FIC_1_ACLK = 0.759"
syn_tsu612 = " FIC_1_AXI4_S_AWADDR[4]->FIC_1_ACLK = 0.765"
syn_tsu613 = " FIC_1_AXI4_S_AWADDR[5]->FIC_1_ACLK = 0.765"
syn_tsu614 = " FIC_1_AXI4_S_AWADDR[6]->FIC_1_ACLK = 0.762"
syn_tsu615 = " FIC_1_AXI4_S_AWADDR[7]->FIC_1_ACLK = 0.76"
syn_tsu616 = " FIC_1_AXI4_S_AWADDR[8]->FIC_1_ACLK = 0.791"
syn_tsu617 = " FIC_1_AXI4_S_AWADDR[9]->FIC_1_ACLK = 0.8"
syn_tsu618 = " FIC_1_AXI4_S_AWBURST[0]->FIC_1_ACLK = 0.764"
syn_tsu619 = " FIC_1_AXI4_S_AWBURST[1]->FIC_1_ACLK = 0.768"
syn_tsu620 = " FIC_1_AXI4_S_AWCACHE[0]->FIC_1_ACLK = 0.755"
syn_tsu621 = " FIC_1_AXI4_S_AWCACHE[1]->FIC_1_ACLK = 0.747"
syn_tsu622 = " FIC_1_AXI4_S_AWCACHE[2]->FIC_1_ACLK = 0.763"
syn_tsu623 = " FIC_1_AXI4_S_AWCACHE[3]->FIC_1_ACLK = 0.778"
syn_tsu624 = " FIC_1_AXI4_S_AWID[0]->FIC_1_ACLK = 0.735"
syn_tsu625 = " FIC_1_AXI4_S_AWID[1]->FIC_1_ACLK = 0.788"
syn_tsu626 = " FIC_1_AXI4_S_AWID[2]->FIC_1_ACLK = 0.752"
syn_tsu627 = " FIC_1_AXI4_S_AWID[3]->FIC_1_ACLK = 0.76"
syn_tsu628 = " FIC_1_AXI4_S_AWLEN[0]->FIC_1_ACLK = 0.772"
syn_tsu629 = " FIC_1_AXI4_S_AWLEN[1]->FIC_1_ACLK = 0.77"
syn_tsu630 = " FIC_1_AXI4_S_AWLEN[2]->FIC_1_ACLK = 0.776"
syn_tsu631 = " FIC_1_AXI4_S_AWLEN[3]->FIC_1_ACLK = 0.801"
syn_tsu632 = " FIC_1_AXI4_S_AWLEN[4]->FIC_1_ACLK = 0.815"
syn_tsu633 = " FIC_1_AXI4_S_AWLEN[5]->FIC_1_ACLK = 0.752"
syn_tsu634 = " FIC_1_AXI4_S_AWLEN[6]->FIC_1_ACLK = 0.743"
syn_tsu635 = " FIC_1_AXI4_S_AWLEN[7]->FIC_1_ACLK = 0.795"
syn_tsu636 = " FIC_1_AXI4_S_AWLOCK->FIC_1_ACLK = 0.772"
syn_tsu637 = " FIC_1_AXI4_S_AWPROT[0]->FIC_1_ACLK = 0.745"
syn_tsu638 = " FIC_1_AXI4_S_AWPROT[1]->FIC_1_ACLK = 0.748"
syn_tsu639 = " FIC_1_AXI4_S_AWPROT[2]->FIC_1_ACLK = 0.729"
syn_tsu640 = " FIC_1_AXI4_S_AWQOS[0]->FIC_1_ACLK = 0.756"
syn_tsu641 = " FIC_1_AXI4_S_AWQOS[1]->FIC_1_ACLK = 0.768"
syn_tsu642 = " FIC_1_AXI4_S_AWQOS[2]->FIC_1_ACLK = 0.713"
syn_tsu643 = " FIC_1_AXI4_S_AWQOS[3]->FIC_1_ACLK = 0.812"
syn_tsu644 = " FIC_1_AXI4_S_AWSIZE[0]->FIC_1_ACLK = 0.753"
syn_tsu645 = " FIC_1_AXI4_S_AWSIZE[1]->FIC_1_ACLK = 0.761"
syn_tsu646 = " FIC_1_AXI4_S_AWSIZE[2]->FIC_1_ACLK = 0.75"
syn_tsu647 = " FIC_1_AXI4_S_AWVALID->FIC_1_ACLK = 0.95"
syn_tsu648 = " FIC_1_AXI4_S_BREADY->FIC_1_ACLK = 0.983"
syn_tsu649 = " FIC_1_AXI4_S_RREADY->FIC_1_ACLK = 1.03"
syn_tsu650 = " FIC_1_AXI4_S_WDATA[0]->FIC_1_ACLK = 1.006"
syn_tsu651 = " FIC_1_AXI4_S_WDATA[10]->FIC_1_ACLK = 0.799"
syn_tsu652 = " FIC_1_AXI4_S_WDATA[11]->FIC_1_ACLK = 0.791"
syn_tsu653 = " FIC_1_AXI4_S_WDATA[12]->FIC_1_ACLK = 0.811"
syn_tsu654 = " FIC_1_AXI4_S_WDATA[13]->FIC_1_ACLK = 0.783"
syn_tsu655 = " FIC_1_AXI4_S_WDATA[14]->FIC_1_ACLK = 0.79"
syn_tsu656 = " FIC_1_AXI4_S_WDATA[15]->FIC_1_ACLK = 0.803"
syn_tsu657 = " FIC_1_AXI4_S_WDATA[16]->FIC_1_ACLK = 0.791"
syn_tsu658 = " FIC_1_AXI4_S_WDATA[17]->FIC_1_ACLK = 0.831"
syn_tsu659 = " FIC_1_AXI4_S_WDATA[18]->FIC_1_ACLK = 0.774"
syn_tsu660 = " FIC_1_AXI4_S_WDATA[19]->FIC_1_ACLK = 0.834"
syn_tsu661 = " FIC_1_AXI4_S_WDATA[1]->FIC_1_ACLK = 0.89"
syn_tsu662 = " FIC_1_AXI4_S_WDATA[20]->FIC_1_ACLK = 0.823"
syn_tsu663 = " FIC_1_AXI4_S_WDATA[21]->FIC_1_ACLK = 0.856"
syn_tsu664 = " FIC_1_AXI4_S_WDATA[22]->FIC_1_ACLK = 0.889"
syn_tsu665 = " FIC_1_AXI4_S_WDATA[23]->FIC_1_ACLK = 0.821"
syn_tsu666 = " FIC_1_AXI4_S_WDATA[24]->FIC_1_ACLK = 0.779"
syn_tsu667 = " FIC_1_AXI4_S_WDATA[25]->FIC_1_ACLK = 0.912"
syn_tsu668 = " FIC_1_AXI4_S_WDATA[26]->FIC_1_ACLK = 0.856"
syn_tsu669 = " FIC_1_AXI4_S_WDATA[27]->FIC_1_ACLK = 0.787"
syn_tsu670 = " FIC_1_AXI4_S_WDATA[28]->FIC_1_ACLK = 0.722"
syn_tsu671 = " FIC_1_AXI4_S_WDATA[29]->FIC_1_ACLK = 0.805"
syn_tsu672 = " FIC_1_AXI4_S_WDATA[2]->FIC_1_ACLK = 0.977"
syn_tsu673 = " FIC_1_AXI4_S_WDATA[30]->FIC_1_ACLK = 0.776"
syn_tsu674 = " FIC_1_AXI4_S_WDATA[31]->FIC_1_ACLK = 0.763"
syn_tsu675 = " FIC_1_AXI4_S_WDATA[32]->FIC_1_ACLK = 0.85"
syn_tsu676 = " FIC_1_AXI4_S_WDATA[33]->FIC_1_ACLK = 0.731"
syn_tsu677 = " FIC_1_AXI4_S_WDATA[34]->FIC_1_ACLK = 0.801"
syn_tsu678 = " FIC_1_AXI4_S_WDATA[35]->FIC_1_ACLK = 0.818"
syn_tsu679 = " FIC_1_AXI4_S_WDATA[36]->FIC_1_ACLK = 0.76"
syn_tsu680 = " FIC_1_AXI4_S_WDATA[37]->FIC_1_ACLK = 0.765"
syn_tsu681 = " FIC_1_AXI4_S_WDATA[38]->FIC_1_ACLK = 0.729"
syn_tsu682 = " FIC_1_AXI4_S_WDATA[39]->FIC_1_ACLK = 0.716"
syn_tsu683 = " FIC_1_AXI4_S_WDATA[3]->FIC_1_ACLK = 0.948"
syn_tsu684 = " FIC_1_AXI4_S_WDATA[40]->FIC_1_ACLK = 0.762"
syn_tsu685 = " FIC_1_AXI4_S_WDATA[41]->FIC_1_ACLK = 0.83"
syn_tsu686 = " FIC_1_AXI4_S_WDATA[42]->FIC_1_ACLK = 0.81"
syn_tsu687 = " FIC_1_AXI4_S_WDATA[43]->FIC_1_ACLK = 0.743"
syn_tsu688 = " FIC_1_AXI4_S_WDATA[44]->FIC_1_ACLK = 0.811"
syn_tsu689 = " FIC_1_AXI4_S_WDATA[45]->FIC_1_ACLK = 0.822"
syn_tsu690 = " FIC_1_AXI4_S_WDATA[46]->FIC_1_ACLK = 0.758"
syn_tsu691 = " FIC_1_AXI4_S_WDATA[47]->FIC_1_ACLK = 0.849"
syn_tsu692 = " FIC_1_AXI4_S_WDATA[48]->FIC_1_ACLK = 0.794"
syn_tsu693 = " FIC_1_AXI4_S_WDATA[49]->FIC_1_ACLK = 0.717"
syn_tsu694 = " FIC_1_AXI4_S_WDATA[4]->FIC_1_ACLK = 0.87"
syn_tsu695 = " FIC_1_AXI4_S_WDATA[50]->FIC_1_ACLK = 0.909"
syn_tsu696 = " FIC_1_AXI4_S_WDATA[51]->FIC_1_ACLK = 0.891"
syn_tsu697 = " FIC_1_AXI4_S_WDATA[52]->FIC_1_ACLK = 0.737"
syn_tsu698 = " FIC_1_AXI4_S_WDATA[53]->FIC_1_ACLK = 0.769"
syn_tsu699 = " FIC_1_AXI4_S_WDATA[54]->FIC_1_ACLK = 0.816"
syn_tsu700 = " FIC_1_AXI4_S_WDATA[55]->FIC_1_ACLK = 0.75"
syn_tsu701 = " FIC_1_AXI4_S_WDATA[56]->FIC_1_ACLK = 0.77"
syn_tsu702 = " FIC_1_AXI4_S_WDATA[57]->FIC_1_ACLK = 0.733"
syn_tsu703 = " FIC_1_AXI4_S_WDATA[58]->FIC_1_ACLK = 0.84"
syn_tsu704 = " FIC_1_AXI4_S_WDATA[59]->FIC_1_ACLK = 0.802"
syn_tsu705 = " FIC_1_AXI4_S_WDATA[5]->FIC_1_ACLK = 0.884"
syn_tsu706 = " FIC_1_AXI4_S_WDATA[60]->FIC_1_ACLK = 0.93"
syn_tsu707 = " FIC_1_AXI4_S_WDATA[61]->FIC_1_ACLK = 0.766"
syn_tsu708 = " FIC_1_AXI4_S_WDATA[62]->FIC_1_ACLK = 0.787"
syn_tsu709 = " FIC_1_AXI4_S_WDATA[63]->FIC_1_ACLK = 0.846"
syn_tsu710 = " FIC_1_AXI4_S_WDATA[6]->FIC_1_ACLK = 0.914"
syn_tsu711 = " FIC_1_AXI4_S_WDATA[7]->FIC_1_ACLK = 0.865"
syn_tsu712 = " FIC_1_AXI4_S_WDATA[8]->FIC_1_ACLK = 0.898"
syn_tsu713 = " FIC_1_AXI4_S_WDATA[9]->FIC_1_ACLK = 0.789"
syn_tsu714 = " FIC_1_AXI4_S_WLAST->FIC_1_ACLK = 0.999"
syn_tsu715 = " FIC_1_AXI4_S_WSTRB[0]->FIC_1_ACLK = 0.972"
syn_tsu716 = " FIC_1_AXI4_S_WSTRB[1]->FIC_1_ACLK = 0.948"
syn_tsu717 = " FIC_1_AXI4_S_WSTRB[2]->FIC_1_ACLK = 1.029"
syn_tsu718 = " FIC_1_AXI4_S_WSTRB[3]->FIC_1_ACLK = 0.979"
syn_tsu719 = " FIC_1_AXI4_S_WSTRB[4]->FIC_1_ACLK = 0.986"
syn_tsu720 = " FIC_1_AXI4_S_WSTRB[5]->FIC_1_ACLK = 0.897"
syn_tsu721 = " FIC_1_AXI4_S_WSTRB[6]->FIC_1_ACLK = 1.005"
syn_tsu722 = " FIC_1_AXI4_S_WSTRB[7]->FIC_1_ACLK = 1.011"
syn_tsu723 = " FIC_1_AXI4_S_WVALID->FIC_1_ACLK = 1.034"
syn_tsu724 = " FIC_2_AXI4_S_ARADDR[0]->FIC_2_ACLK = 0.768"
syn_tsu725 = " FIC_2_AXI4_S_ARADDR[10]->FIC_2_ACLK = 0.83"
syn_tsu726 = " FIC_2_AXI4_S_ARADDR[11]->FIC_2_ACLK = 0.847"
syn_tsu727 = " FIC_2_AXI4_S_ARADDR[12]->FIC_2_ACLK = 0.835"
syn_tsu728 = " FIC_2_AXI4_S_ARADDR[13]->FIC_2_ACLK = 0.852"
syn_tsu729 = " FIC_2_AXI4_S_ARADDR[14]->FIC_2_ACLK = 0.818"
syn_tsu730 = " FIC_2_AXI4_S_ARADDR[15]->FIC_2_ACLK = 0.819"
syn_tsu731 = " FIC_2_AXI4_S_ARADDR[16]->FIC_2_ACLK = 0.82"
syn_tsu732 = " FIC_2_AXI4_S_ARADDR[17]->FIC_2_ACLK = 0.833"
syn_tsu733 = " FIC_2_AXI4_S_ARADDR[18]->FIC_2_ACLK = 0.879"
syn_tsu734 = " FIC_2_AXI4_S_ARADDR[19]->FIC_2_ACLK = 0.848"
syn_tsu735 = " FIC_2_AXI4_S_ARADDR[1]->FIC_2_ACLK = 0.769"
syn_tsu736 = " FIC_2_AXI4_S_ARADDR[20]->FIC_2_ACLK = 0.87"
syn_tsu737 = " FIC_2_AXI4_S_ARADDR[21]->FIC_2_ACLK = 0.867"
syn_tsu738 = " FIC_2_AXI4_S_ARADDR[22]->FIC_2_ACLK = 0.84"
syn_tsu739 = " FIC_2_AXI4_S_ARADDR[23]->FIC_2_ACLK = 0.861"
syn_tsu740 = " FIC_2_AXI4_S_ARADDR[24]->FIC_2_ACLK = 0.838"
syn_tsu741 = " FIC_2_AXI4_S_ARADDR[25]->FIC_2_ACLK = 0.865"
syn_tsu742 = " FIC_2_AXI4_S_ARADDR[26]->FIC_2_ACLK = 0.841"
syn_tsu743 = " FIC_2_AXI4_S_ARADDR[27]->FIC_2_ACLK = 0.86"
syn_tsu744 = " FIC_2_AXI4_S_ARADDR[28]->FIC_2_ACLK = 0.837"
syn_tsu745 = " FIC_2_AXI4_S_ARADDR[29]->FIC_2_ACLK = 0.821"
syn_tsu746 = " FIC_2_AXI4_S_ARADDR[2]->FIC_2_ACLK = 0.803"
syn_tsu747 = " FIC_2_AXI4_S_ARADDR[30]->FIC_2_ACLK = 0.801"
syn_tsu748 = " FIC_2_AXI4_S_ARADDR[31]->FIC_2_ACLK = 0.807"
syn_tsu749 = " FIC_2_AXI4_S_ARADDR[32]->FIC_2_ACLK = 0.817"
syn_tsu750 = " FIC_2_AXI4_S_ARADDR[33]->FIC_2_ACLK = 0.821"
syn_tsu751 = " FIC_2_AXI4_S_ARADDR[34]->FIC_2_ACLK = 0.836"
syn_tsu752 = " FIC_2_AXI4_S_ARADDR[35]->FIC_2_ACLK = 0.838"
syn_tsu753 = " FIC_2_AXI4_S_ARADDR[36]->FIC_2_ACLK = 0.811"
syn_tsu754 = " FIC_2_AXI4_S_ARADDR[37]->FIC_2_ACLK = 0.818"
syn_tsu755 = " FIC_2_AXI4_S_ARADDR[3]->FIC_2_ACLK = 0.817"
syn_tsu756 = " FIC_2_AXI4_S_ARADDR[4]->FIC_2_ACLK = 0.803"
syn_tsu757 = " FIC_2_AXI4_S_ARADDR[5]->FIC_2_ACLK = 0.79"
syn_tsu758 = " FIC_2_AXI4_S_ARADDR[6]->FIC_2_ACLK = 0.77"
syn_tsu759 = " FIC_2_AXI4_S_ARADDR[7]->FIC_2_ACLK = 0.786"
syn_tsu760 = " FIC_2_AXI4_S_ARADDR[8]->FIC_2_ACLK = 0.796"
syn_tsu761 = " FIC_2_AXI4_S_ARADDR[9]->FIC_2_ACLK = 0.818"
syn_tsu762 = " FIC_2_AXI4_S_ARBURST[0]->FIC_2_ACLK = 0.808"
syn_tsu763 = " FIC_2_AXI4_S_ARBURST[1]->FIC_2_ACLK = 0.797"
syn_tsu764 = " FIC_2_AXI4_S_ARID[0]->FIC_2_ACLK = 0.84"
syn_tsu765 = " FIC_2_AXI4_S_ARID[1]->FIC_2_ACLK = 0.814"
syn_tsu766 = " FIC_2_AXI4_S_ARID[2]->FIC_2_ACLK = 0.824"
syn_tsu767 = " FIC_2_AXI4_S_ARID[3]->FIC_2_ACLK = 0.821"
syn_tsu768 = " FIC_2_AXI4_S_ARLEN[0]->FIC_2_ACLK = 0.772"
syn_tsu769 = " FIC_2_AXI4_S_ARLEN[1]->FIC_2_ACLK = 0.804"
syn_tsu770 = " FIC_2_AXI4_S_ARLEN[2]->FIC_2_ACLK = 0.762"
syn_tsu771 = " FIC_2_AXI4_S_ARLEN[3]->FIC_2_ACLK = 0.786"
syn_tsu772 = " FIC_2_AXI4_S_ARLEN[4]->FIC_2_ACLK = 0.796"
syn_tsu773 = " FIC_2_AXI4_S_ARLEN[5]->FIC_2_ACLK = 0.789"
syn_tsu774 = " FIC_2_AXI4_S_ARLEN[6]->FIC_2_ACLK = 0.874"
syn_tsu775 = " FIC_2_AXI4_S_ARLEN[7]->FIC_2_ACLK = 0.8"
syn_tsu776 = " FIC_2_AXI4_S_ARLOCK->FIC_2_ACLK = 0.823"
syn_tsu777 = " FIC_2_AXI4_S_ARPROT[0]->FIC_2_ACLK = 0.808"
syn_tsu778 = " FIC_2_AXI4_S_ARPROT[1]->FIC_2_ACLK = 0.799"
syn_tsu779 = " FIC_2_AXI4_S_ARPROT[2]->FIC_2_ACLK = 0.789"
syn_tsu780 = " FIC_2_AXI4_S_ARQOS[0]->FIC_2_ACLK = 0.793"
syn_tsu781 = " FIC_2_AXI4_S_ARQOS[1]->FIC_2_ACLK = 0.791"
syn_tsu782 = " FIC_2_AXI4_S_ARQOS[2]->FIC_2_ACLK = 0.778"
syn_tsu783 = " FIC_2_AXI4_S_ARQOS[3]->FIC_2_ACLK = 0.779"
syn_tsu784 = " FIC_2_AXI4_S_ARSIZE[0]->FIC_2_ACLK = 0.838"
syn_tsu785 = " FIC_2_AXI4_S_ARSIZE[1]->FIC_2_ACLK = 0.819"
syn_tsu786 = " FIC_2_AXI4_S_ARSIZE[2]->FIC_2_ACLK = 0.796"
syn_tsu787 = " FIC_2_AXI4_S_ARVALID->FIC_2_ACLK = 1.088"
syn_tsu788 = " FIC_2_AXI4_S_AWADDR[0]->FIC_2_ACLK = 0.873"
syn_tsu789 = " FIC_2_AXI4_S_AWADDR[10]->FIC_2_ACLK = 0.829"
syn_tsu790 = " FIC_2_AXI4_S_AWADDR[11]->FIC_2_ACLK = 0.878"
syn_tsu791 = " FIC_2_AXI4_S_AWADDR[12]->FIC_2_ACLK = 0.846"
syn_tsu792 = " FIC_2_AXI4_S_AWADDR[13]->FIC_2_ACLK = 0.863"
syn_tsu793 = " FIC_2_AXI4_S_AWADDR[14]->FIC_2_ACLK = 0.822"
syn_tsu794 = " FIC_2_AXI4_S_AWADDR[15]->FIC_2_ACLK = 0.779"
syn_tsu795 = " FIC_2_AXI4_S_AWADDR[16]->FIC_2_ACLK = 0.826"
syn_tsu796 = " FIC_2_AXI4_S_AWADDR[17]->FIC_2_ACLK = 0.804"
syn_tsu797 = " FIC_2_AXI4_S_AWADDR[18]->FIC_2_ACLK = 0.824"
syn_tsu798 = " FIC_2_AXI4_S_AWADDR[19]->FIC_2_ACLK = 0.815"
syn_tsu799 = " FIC_2_AXI4_S_AWADDR[1]->FIC_2_ACLK = 0.861"
syn_tsu800 = " FIC_2_AXI4_S_AWADDR[20]->FIC_2_ACLK = 0.797"
syn_tsu801 = " FIC_2_AXI4_S_AWADDR[21]->FIC_2_ACLK = 0.822"
syn_tsu802 = " FIC_2_AXI4_S_AWADDR[22]->FIC_2_ACLK = 0.789"
syn_tsu803 = " FIC_2_AXI4_S_AWADDR[23]->FIC_2_ACLK = 0.777"
syn_tsu804 = " FIC_2_AXI4_S_AWADDR[24]->FIC_2_ACLK = 0.768"
syn_tsu805 = " FIC_2_AXI4_S_AWADDR[25]->FIC_2_ACLK = 0.76"
syn_tsu806 = " FIC_2_AXI4_S_AWADDR[26]->FIC_2_ACLK = 0.774"
syn_tsu807 = " FIC_2_AXI4_S_AWADDR[27]->FIC_2_ACLK = 0.818"
syn_tsu808 = " FIC_2_AXI4_S_AWADDR[28]->FIC_2_ACLK = 0.79"
syn_tsu809 = " FIC_2_AXI4_S_AWADDR[29]->FIC_2_ACLK = 0.789"
syn_tsu810 = " FIC_2_AXI4_S_AWADDR[2]->FIC_2_ACLK = 0.909"
syn_tsu811 = " FIC_2_AXI4_S_AWADDR[30]->FIC_2_ACLK = 0.797"
syn_tsu812 = " FIC_2_AXI4_S_AWADDR[31]->FIC_2_ACLK = 0.791"
syn_tsu813 = " FIC_2_AXI4_S_AWADDR[32]->FIC_2_ACLK = 0.801"
syn_tsu814 = " FIC_2_AXI4_S_AWADDR[33]->FIC_2_ACLK = 0.816"
syn_tsu815 = " FIC_2_AXI4_S_AWADDR[34]->FIC_2_ACLK = 0.811"
syn_tsu816 = " FIC_2_AXI4_S_AWADDR[35]->FIC_2_ACLK = 0.817"
syn_tsu817 = " FIC_2_AXI4_S_AWADDR[36]->FIC_2_ACLK = 0.807"
syn_tsu818 = " FIC_2_AXI4_S_AWADDR[37]->FIC_2_ACLK = 0.789"
syn_tsu819 = " FIC_2_AXI4_S_AWADDR[3]->FIC_2_ACLK = 0.909"
syn_tsu820 = " FIC_2_AXI4_S_AWADDR[4]->FIC_2_ACLK = 0.87"
syn_tsu821 = " FIC_2_AXI4_S_AWADDR[5]->FIC_2_ACLK = 0.921"
syn_tsu822 = " FIC_2_AXI4_S_AWADDR[6]->FIC_2_ACLK = 0.88"
syn_tsu823 = " FIC_2_AXI4_S_AWADDR[7]->FIC_2_ACLK = 0.859"
syn_tsu824 = " FIC_2_AXI4_S_AWADDR[8]->FIC_2_ACLK = 0.853"
syn_tsu825 = " FIC_2_AXI4_S_AWADDR[9]->FIC_2_ACLK = 0.827"
syn_tsu826 = " FIC_2_AXI4_S_AWBURST[0]->FIC_2_ACLK = 0.885"
syn_tsu827 = " FIC_2_AXI4_S_AWBURST[1]->FIC_2_ACLK = 0.938"
syn_tsu828 = " FIC_2_AXI4_S_AWID[0]->FIC_2_ACLK = 0.852"
syn_tsu829 = " FIC_2_AXI4_S_AWID[1]->FIC_2_ACLK = 0.819"
syn_tsu830 = " FIC_2_AXI4_S_AWID[2]->FIC_2_ACLK = 0.834"
syn_tsu831 = " FIC_2_AXI4_S_AWID[3]->FIC_2_ACLK = 0.852"
syn_tsu832 = " FIC_2_AXI4_S_AWLEN[0]->FIC_2_ACLK = 0.885"
syn_tsu833 = " FIC_2_AXI4_S_AWLEN[1]->FIC_2_ACLK = 0.979"
syn_tsu834 = " FIC_2_AXI4_S_AWLEN[2]->FIC_2_ACLK = 1.033"
syn_tsu835 = " FIC_2_AXI4_S_AWLEN[3]->FIC_2_ACLK = 1.031"
syn_tsu836 = " FIC_2_AXI4_S_AWLEN[4]->FIC_2_ACLK = 0.839"
syn_tsu837 = " FIC_2_AXI4_S_AWLEN[5]->FIC_2_ACLK = 0.925"
syn_tsu838 = " FIC_2_AXI4_S_AWLEN[6]->FIC_2_ACLK = 0.884"
syn_tsu839 = " FIC_2_AXI4_S_AWLEN[7]->FIC_2_ACLK = 0.877"
syn_tsu840 = " FIC_2_AXI4_S_AWLOCK->FIC_2_ACLK = 0.993"
syn_tsu841 = " FIC_2_AXI4_S_AWPROT[0]->FIC_2_ACLK = 1.013"
syn_tsu842 = " FIC_2_AXI4_S_AWPROT[1]->FIC_2_ACLK = 1.012"
syn_tsu843 = " FIC_2_AXI4_S_AWPROT[2]->FIC_2_ACLK = 1.002"
syn_tsu844 = " FIC_2_AXI4_S_AWQOS[0]->FIC_2_ACLK = 1.004"
syn_tsu845 = " FIC_2_AXI4_S_AWQOS[1]->FIC_2_ACLK = 1.004"
syn_tsu846 = " FIC_2_AXI4_S_AWQOS[2]->FIC_2_ACLK = 1.009"
syn_tsu847 = " FIC_2_AXI4_S_AWQOS[3]->FIC_2_ACLK = 0.987"
syn_tsu848 = " FIC_2_AXI4_S_AWSIZE[0]->FIC_2_ACLK = 0.974"
syn_tsu849 = " FIC_2_AXI4_S_AWSIZE[1]->FIC_2_ACLK = 0.983"
syn_tsu850 = " FIC_2_AXI4_S_AWSIZE[2]->FIC_2_ACLK = 1.041"
syn_tsu851 = " FIC_2_AXI4_S_AWVALID->FIC_2_ACLK = 1.033"
syn_tsu852 = " FIC_2_AXI4_S_BREADY->FIC_2_ACLK = 1.046"
syn_tsu853 = " FIC_2_AXI4_S_RREADY->FIC_2_ACLK = 1.027"
syn_tsu854 = " FIC_2_AXI4_S_WDATA[0]->FIC_2_ACLK = 0.963"
syn_tsu855 = " FIC_2_AXI4_S_WDATA[10]->FIC_2_ACLK = 0.951"
syn_tsu856 = " FIC_2_AXI4_S_WDATA[11]->FIC_2_ACLK = 0.982"
syn_tsu857 = " FIC_2_AXI4_S_WDATA[12]->FIC_2_ACLK = 0.959"
syn_tsu858 = " FIC_2_AXI4_S_WDATA[13]->FIC_2_ACLK = 0.884"
syn_tsu859 = " FIC_2_AXI4_S_WDATA[14]->FIC_2_ACLK = 0.975"
syn_tsu860 = " FIC_2_AXI4_S_WDATA[15]->FIC_2_ACLK = 0.997"
syn_tsu861 = " FIC_2_AXI4_S_WDATA[16]->FIC_2_ACLK = 0.986"
syn_tsu862 = " FIC_2_AXI4_S_WDATA[17]->FIC_2_ACLK = 0.988"
syn_tsu863 = " FIC_2_AXI4_S_WDATA[18]->FIC_2_ACLK = 0.985"
syn_tsu864 = " FIC_2_AXI4_S_WDATA[19]->FIC_2_ACLK = 0.891"
syn_tsu865 = " FIC_2_AXI4_S_WDATA[1]->FIC_2_ACLK = 0.998"
syn_tsu866 = " FIC_2_AXI4_S_WDATA[20]->FIC_2_ACLK = 0.981"
syn_tsu867 = " FIC_2_AXI4_S_WDATA[21]->FIC_2_ACLK = 1.078"
syn_tsu868 = " FIC_2_AXI4_S_WDATA[22]->FIC_2_ACLK = 0.982"
syn_tsu869 = " FIC_2_AXI4_S_WDATA[23]->FIC_2_ACLK = 0.983"
syn_tsu870 = " FIC_2_AXI4_S_WDATA[24]->FIC_2_ACLK = 1.001"
syn_tsu871 = " FIC_2_AXI4_S_WDATA[25]->FIC_2_ACLK = 0.994"
syn_tsu872 = " FIC_2_AXI4_S_WDATA[26]->FIC_2_ACLK = 1.018"
syn_tsu873 = " FIC_2_AXI4_S_WDATA[27]->FIC_2_ACLK = 0.97"
syn_tsu874 = " FIC_2_AXI4_S_WDATA[28]->FIC_2_ACLK = 0.948"
syn_tsu875 = " FIC_2_AXI4_S_WDATA[29]->FIC_2_ACLK = 0.966"
syn_tsu876 = " FIC_2_AXI4_S_WDATA[2]->FIC_2_ACLK = 0.989"
syn_tsu877 = " FIC_2_AXI4_S_WDATA[30]->FIC_2_ACLK = 0.901"
syn_tsu878 = " FIC_2_AXI4_S_WDATA[31]->FIC_2_ACLK = 0.972"
syn_tsu879 = " FIC_2_AXI4_S_WDATA[32]->FIC_2_ACLK = 1.038"
syn_tsu880 = " FIC_2_AXI4_S_WDATA[33]->FIC_2_ACLK = 0.937"
syn_tsu881 = " FIC_2_AXI4_S_WDATA[34]->FIC_2_ACLK = 1.016"
syn_tsu882 = " FIC_2_AXI4_S_WDATA[35]->FIC_2_ACLK = 0.985"
syn_tsu883 = " FIC_2_AXI4_S_WDATA[36]->FIC_2_ACLK = 1.056"
syn_tsu884 = " FIC_2_AXI4_S_WDATA[37]->FIC_2_ACLK = 0.959"
syn_tsu885 = " FIC_2_AXI4_S_WDATA[38]->FIC_2_ACLK = 1.011"
syn_tsu886 = " FIC_2_AXI4_S_WDATA[39]->FIC_2_ACLK = 1.068"
syn_tsu887 = " FIC_2_AXI4_S_WDATA[3]->FIC_2_ACLK = 0.996"
syn_tsu888 = " FIC_2_AXI4_S_WDATA[40]->FIC_2_ACLK = 0.99"
syn_tsu889 = " FIC_2_AXI4_S_WDATA[41]->FIC_2_ACLK = 1.063"
syn_tsu890 = " FIC_2_AXI4_S_WDATA[42]->FIC_2_ACLK = 0.98"
syn_tsu891 = " FIC_2_AXI4_S_WDATA[43]->FIC_2_ACLK = 1.013"
syn_tsu892 = " FIC_2_AXI4_S_WDATA[44]->FIC_2_ACLK = 0.965"
syn_tsu893 = " FIC_2_AXI4_S_WDATA[45]->FIC_2_ACLK = 1.011"
syn_tsu894 = " FIC_2_AXI4_S_WDATA[46]->FIC_2_ACLK = 0.983"
syn_tsu895 = " FIC_2_AXI4_S_WDATA[47]->FIC_2_ACLK = 1.032"
syn_tsu896 = " FIC_2_AXI4_S_WDATA[48]->FIC_2_ACLK = 0.996"
syn_tsu897 = " FIC_2_AXI4_S_WDATA[49]->FIC_2_ACLK = 0.975"
syn_tsu898 = " FIC_2_AXI4_S_WDATA[4]->FIC_2_ACLK = 0.951"
syn_tsu899 = " FIC_2_AXI4_S_WDATA[50]->FIC_2_ACLK = 1.046"
syn_tsu900 = " FIC_2_AXI4_S_WDATA[51]->FIC_2_ACLK = 0.883"
syn_tsu901 = " FIC_2_AXI4_S_WDATA[52]->FIC_2_ACLK = 0.997"
syn_tsu902 = " FIC_2_AXI4_S_WDATA[53]->FIC_2_ACLK = 0.919"
syn_tsu903 = " FIC_2_AXI4_S_WDATA[54]->FIC_2_ACLK = 0.979"
syn_tsu904 = " FIC_2_AXI4_S_WDATA[55]->FIC_2_ACLK = 0.823"
syn_tsu905 = " FIC_2_AXI4_S_WDATA[56]->FIC_2_ACLK = 0.925"
syn_tsu906 = " FIC_2_AXI4_S_WDATA[57]->FIC_2_ACLK = 0.928"
syn_tsu907 = " FIC_2_AXI4_S_WDATA[58]->FIC_2_ACLK = 0.91"
syn_tsu908 = " FIC_2_AXI4_S_WDATA[59]->FIC_2_ACLK = 0.98"
syn_tsu909 = " FIC_2_AXI4_S_WDATA[5]->FIC_2_ACLK = 1.006"
syn_tsu910 = " FIC_2_AXI4_S_WDATA[60]->FIC_2_ACLK = 0.946"
syn_tsu911 = " FIC_2_AXI4_S_WDATA[61]->FIC_2_ACLK = 0.986"
syn_tsu912 = " FIC_2_AXI4_S_WDATA[62]->FIC_2_ACLK = 0.861"
syn_tsu913 = " FIC_2_AXI4_S_WDATA[63]->FIC_2_ACLK = 1.033"
syn_tsu914 = " FIC_2_AXI4_S_WDATA[6]->FIC_2_ACLK = 0.964"
syn_tsu915 = " FIC_2_AXI4_S_WDATA[7]->FIC_2_ACLK = 1.063"
syn_tsu916 = " FIC_2_AXI4_S_WDATA[8]->FIC_2_ACLK = 0.966"
syn_tsu917 = " FIC_2_AXI4_S_WDATA[9]->FIC_2_ACLK = 0.94"
syn_tsu918 = " FIC_2_AXI4_S_WLAST->FIC_2_ACLK = 0.979"
syn_tsu919 = " FIC_2_AXI4_S_WSTRB[0]->FIC_2_ACLK = 1.043"
syn_tsu920 = " FIC_2_AXI4_S_WSTRB[1]->FIC_2_ACLK = 0.98"
syn_tsu921 = " FIC_2_AXI4_S_WSTRB[2]->FIC_2_ACLK = 0.97"
syn_tsu922 = " FIC_2_AXI4_S_WSTRB[3]->FIC_2_ACLK = 0.978"
syn_tsu923 = " FIC_2_AXI4_S_WSTRB[4]->FIC_2_ACLK = 1.001"
syn_tsu924 = " FIC_2_AXI4_S_WSTRB[5]->FIC_2_ACLK = 0.983"
syn_tsu925 = " FIC_2_AXI4_S_WSTRB[6]->FIC_2_ACLK = 0.976"
syn_tsu926 = " FIC_2_AXI4_S_WSTRB[7]->FIC_2_ACLK = 0.992"
syn_tsu927 = " FIC_2_AXI4_S_WVALID->FIC_2_ACLK = 1.064"
syn_tsu928 = " FIC_3_APB_M_PRDATA[0]->FIC_3_PCLK = 0"
syn_tsu929 = " FIC_3_APB_M_PRDATA[10]->FIC_3_PCLK = 0"
syn_tsu930 = " FIC_3_APB_M_PRDATA[11]->FIC_3_PCLK = 0"
syn_tsu931 = " FIC_3_APB_M_PRDATA[12]->FIC_3_PCLK = 0"
syn_tsu932 = " FIC_3_APB_M_PRDATA[13]->FIC_3_PCLK = 0"
syn_tsu933 = " FIC_3_APB_M_PRDATA[14]->FIC_3_PCLK = 0"
syn_tsu934 = " FIC_3_APB_M_PRDATA[15]->FIC_3_PCLK = 0"
syn_tsu935 = " FIC_3_APB_M_PRDATA[16]->FIC_3_PCLK = 0"
syn_tsu936 = " FIC_3_APB_M_PRDATA[17]->FIC_3_PCLK = 0"
syn_tsu937 = " FIC_3_APB_M_PRDATA[18]->FIC_3_PCLK = 0"
syn_tsu938 = " FIC_3_APB_M_PRDATA[19]->FIC_3_PCLK = 0"
syn_tsu939 = " FIC_3_APB_M_PRDATA[1]->FIC_3_PCLK = 0"
syn_tsu940 = " FIC_3_APB_M_PRDATA[20]->FIC_3_PCLK = 0"
syn_tsu941 = " FIC_3_APB_M_PRDATA[21]->FIC_3_PCLK = 0"
syn_tsu942 = " FIC_3_APB_M_PRDATA[22]->FIC_3_PCLK = 0"
syn_tsu943 = " FIC_3_APB_M_PRDATA[23]->FIC_3_PCLK = 0"
syn_tsu944 = " FIC_3_APB_M_PRDATA[24]->FIC_3_PCLK = 0"
syn_tsu945 = " FIC_3_APB_M_PRDATA[25]->FIC_3_PCLK = 0"
syn_tsu946 = " FIC_3_APB_M_PRDATA[26]->FIC_3_PCLK = 0"
syn_tsu947 = " FIC_3_APB_M_PRDATA[27]->FIC_3_PCLK = 0"
syn_tsu948 = " FIC_3_APB_M_PRDATA[28]->FIC_3_PCLK = 0"
syn_tsu949 = " FIC_3_APB_M_PRDATA[29]->FIC_3_PCLK = 0"
syn_tsu950 = " FIC_3_APB_M_PRDATA[2]->FIC_3_PCLK = 0"
syn_tsu951 = " FIC_3_APB_M_PRDATA[30]->FIC_3_PCLK = 0"
syn_tsu952 = " FIC_3_APB_M_PRDATA[31]->FIC_3_PCLK = 0"
syn_tsu953 = " FIC_3_APB_M_PRDATA[3]->FIC_3_PCLK = 0"
syn_tsu954 = " FIC_3_APB_M_PRDATA[4]->FIC_3_PCLK = 0"
syn_tsu955 = " FIC_3_APB_M_PRDATA[5]->FIC_3_PCLK = 0"
syn_tsu956 = " FIC_3_APB_M_PRDATA[6]->FIC_3_PCLK = 0"
syn_tsu957 = " FIC_3_APB_M_PRDATA[7]->FIC_3_PCLK = 0"
syn_tsu958 = " FIC_3_APB_M_PRDATA[8]->FIC_3_PCLK = 0"
syn_tsu959 = " FIC_3_APB_M_PRDATA[9]->FIC_3_PCLK = 0"
syn_tsu960 = " FIC_3_APB_M_PREADY->FIC_3_PCLK = 0"
syn_tsu961 = " FIC_3_APB_M_PSLVERR->FIC_3_PCLK = 0"
syn_tsu962 = " JTAG_TDI_F2M->JTAG_TCK_F2M = 0.894"
syn_tsu963 = " JTAG_TMS_F2M->JTAG_TCK_F2M = 1.759"
syn_tsu964 = " MAC_0_GMII_MII_RXD_F2M[0]->MAC_0_GMII_MII_RX_CLK_F2M = 2.944"
syn_tsu965 = " MAC_0_GMII_MII_RXD_F2M[1]->MAC_0_GMII_MII_RX_CLK_F2M = 2.958"
syn_tsu966 = " MAC_0_GMII_MII_RXD_F2M[2]->MAC_0_GMII_MII_RX_CLK_F2M = 2.928"
syn_tsu967 = " MAC_0_GMII_MII_RXD_F2M[3]->MAC_0_GMII_MII_RX_CLK_F2M = 2.968"
syn_tsu968 = " MAC_0_GMII_MII_RXD_F2M[4]->MAC_0_GMII_MII_RX_CLK_F2M = 2.958"
syn_tsu969 = " MAC_0_GMII_MII_RXD_F2M[5]->MAC_0_GMII_MII_RX_CLK_F2M = 2.995"
syn_tsu970 = " MAC_0_GMII_MII_RXD_F2M[6]->MAC_0_GMII_MII_RX_CLK_F2M = 2.96"
syn_tsu971 = " MAC_0_GMII_MII_RXD_F2M[7]->MAC_0_GMII_MII_RX_CLK_F2M = 3.001"
syn_tsu972 = " MAC_0_GMII_MII_RX_DV_F2M->MAC_0_GMII_MII_RX_CLK_F2M = 2.919"
syn_tsu973 = " MAC_0_GMII_MII_RX_ER_F2M->MAC_0_GMII_MII_RX_CLK_F2M = 2.97"
syn_tsu974 = " MAC_1_GMII_MII_RXD_F2M[0]->MAC_1_GMII_MII_RX_CLK_F2M = 2.811"
syn_tsu975 = " MAC_1_GMII_MII_RXD_F2M[1]->MAC_1_GMII_MII_RX_CLK_F2M = 2.783"
syn_tsu976 = " MAC_1_GMII_MII_RXD_F2M[2]->MAC_1_GMII_MII_RX_CLK_F2M = 2.878"
syn_tsu977 = " MAC_1_GMII_MII_RXD_F2M[3]->MAC_1_GMII_MII_RX_CLK_F2M = 2.79"
syn_tsu978 = " MAC_1_GMII_MII_RXD_F2M[4]->MAC_1_GMII_MII_RX_CLK_F2M = 2.823"
syn_tsu979 = " MAC_1_GMII_MII_RXD_F2M[5]->MAC_1_GMII_MII_RX_CLK_F2M = 2.885"
syn_tsu980 = " MAC_1_GMII_MII_RXD_F2M[6]->MAC_1_GMII_MII_RX_CLK_F2M = 2.834"
syn_tsu981 = " MAC_1_GMII_MII_RXD_F2M[7]->MAC_1_GMII_MII_RX_CLK_F2M = 2.802"
syn_tsu982 = " MAC_1_GMII_MII_RX_DV_F2M->MAC_1_GMII_MII_RX_CLK_F2M = 2.76"
syn_tsu983 = " MAC_1_GMII_MII_RX_ER_F2M->MAC_1_GMII_MII_RX_CLK_F2M = 2.809"
syn_tsu984 = " USOC_TRACE_DATA_F2M[0]->USOC_TRACE_CLOCK_F2M = 0.679"
syn_tsu985 = " USOC_TRACE_DATA_F2M[10]->USOC_TRACE_CLOCK_F2M = 0.812"
syn_tsu986 = " USOC_TRACE_DATA_F2M[11]->USOC_TRACE_CLOCK_F2M = 0.718"
syn_tsu987 = " USOC_TRACE_DATA_F2M[12]->USOC_TRACE_CLOCK_F2M = 0.772"
syn_tsu988 = " USOC_TRACE_DATA_F2M[13]->USOC_TRACE_CLOCK_F2M = 0.777"
syn_tsu989 = " USOC_TRACE_DATA_F2M[14]->USOC_TRACE_CLOCK_F2M = 0.791"
syn_tsu990 = " USOC_TRACE_DATA_F2M[15]->USOC_TRACE_CLOCK_F2M = 0.697"
syn_tsu991 = " USOC_TRACE_DATA_F2M[16]->USOC_TRACE_CLOCK_F2M = 0.7"
syn_tsu992 = " USOC_TRACE_DATA_F2M[17]->USOC_TRACE_CLOCK_F2M = 0.797"
syn_tsu993 = " USOC_TRACE_DATA_F2M[18]->USOC_TRACE_CLOCK_F2M = 0.785"
syn_tsu994 = " USOC_TRACE_DATA_F2M[19]->USOC_TRACE_CLOCK_F2M = 0.793"
syn_tsu995 = " USOC_TRACE_DATA_F2M[1]->USOC_TRACE_CLOCK_F2M = 0.739"
syn_tsu996 = " USOC_TRACE_DATA_F2M[20]->USOC_TRACE_CLOCK_F2M = 0.807"
syn_tsu997 = " USOC_TRACE_DATA_F2M[21]->USOC_TRACE_CLOCK_F2M = 0.708"
syn_tsu998 = " USOC_TRACE_DATA_F2M[22]->USOC_TRACE_CLOCK_F2M = 0.781"
syn_tsu999 = " USOC_TRACE_DATA_F2M[23]->USOC_TRACE_CLOCK_F2M = 0.732"
syn_tsu1000 = " USOC_TRACE_DATA_F2M[24]->USOC_TRACE_CLOCK_F2M = 0.679"
syn_tsu1001 = " USOC_TRACE_DATA_F2M[25]->USOC_TRACE_CLOCK_F2M = 0.656"
syn_tsu1002 = " USOC_TRACE_DATA_F2M[26]->USOC_TRACE_CLOCK_F2M = 0.801"
syn_tsu1003 = " USOC_TRACE_DATA_F2M[27]->USOC_TRACE_CLOCK_F2M = 0.791"
syn_tsu1004 = " USOC_TRACE_DATA_F2M[28]->USOC_TRACE_CLOCK_F2M = 0.764"
syn_tsu1005 = " USOC_TRACE_DATA_F2M[29]->USOC_TRACE_CLOCK_F2M = 0.692"
syn_tsu1006 = " USOC_TRACE_DATA_F2M[2]->USOC_TRACE_CLOCK_F2M = 0.779"
syn_tsu1007 = " USOC_TRACE_DATA_F2M[30]->USOC_TRACE_CLOCK_F2M = 0.727"
syn_tsu1008 = " USOC_TRACE_DATA_F2M[31]->USOC_TRACE_CLOCK_F2M = 0.726"
syn_tsu1009 = " USOC_TRACE_DATA_F2M[32]->USOC_TRACE_CLOCK_F2M = 0.66"
syn_tsu1010 = " USOC_TRACE_DATA_F2M[33]->USOC_TRACE_CLOCK_F2M = 0.753"
syn_tsu1011 = " USOC_TRACE_DATA_F2M[34]->USOC_TRACE_CLOCK_F2M = 0.741"
syn_tsu1012 = " USOC_TRACE_DATA_F2M[35]->USOC_TRACE_CLOCK_F2M = 0.709"
syn_tsu1013 = " USOC_TRACE_DATA_F2M[36]->USOC_TRACE_CLOCK_F2M = 0.655"
syn_tsu1014 = " USOC_TRACE_DATA_F2M[37]->USOC_TRACE_CLOCK_F2M = 0.723"
syn_tsu1015 = " USOC_TRACE_DATA_F2M[38]->USOC_TRACE_CLOCK_F2M = 0.702"
syn_tsu1016 = " USOC_TRACE_DATA_F2M[39]->USOC_TRACE_CLOCK_F2M = 0.717"
syn_tsu1017 = " USOC_TRACE_DATA_F2M[3]->USOC_TRACE_CLOCK_F2M = 0.718"
syn_tsu1018 = " USOC_TRACE_DATA_F2M[4]->USOC_TRACE_CLOCK_F2M = 0.694"
syn_tsu1019 = " USOC_TRACE_DATA_F2M[5]->USOC_TRACE_CLOCK_F2M = 0.714"
syn_tsu1020 = " USOC_TRACE_DATA_F2M[6]->USOC_TRACE_CLOCK_F2M = 0.683"
syn_tsu1021 = " USOC_TRACE_DATA_F2M[7]->USOC_TRACE_CLOCK_F2M = 0.702"
syn_tsu1022 = " USOC_TRACE_DATA_F2M[8]->USOC_TRACE_CLOCK_F2M = 0.75"
syn_tsu1023 = " USOC_TRACE_DATA_F2M[9]->USOC_TRACE_CLOCK_F2M = 0.733"
syn_tsu1024 = " USOC_TRACE_VALID_F2M->USOC_TRACE_CLOCK_F2M = 0.702"
syn_tco0 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[0] = 2.673"
syn_tco1 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[10] = 2.625"
syn_tco2 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[11] = 2.567"
syn_tco3 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[12] = 2.669"
syn_tco4 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[13] = 2.544"
syn_tco5 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[14] = 2.614"
syn_tco6 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[15] = 2.703"
syn_tco7 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[16] = 2.674"
syn_tco8 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[17] = 2.629"
syn_tco9 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[18] = 2.627"
syn_tco10 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[19] = 2.604"
syn_tco11 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[1] = 2.597"
syn_tco12 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[20] = 2.593"
syn_tco13 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[21] = 2.542"
syn_tco14 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[22] = 2.586"
syn_tco15 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[23] = 2.584"
syn_tco16 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[24] = 2.580"
syn_tco17 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[25] = 2.537"
syn_tco18 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[26] = 2.522"
syn_tco19 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[27] = 2.630"
syn_tco20 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[28] = 2.629"
syn_tco21 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[29] = 2.614"
syn_tco22 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[2] = 2.637"
syn_tco23 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[30] = 2.625"
syn_tco24 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[31] = 2.616"
syn_tco25 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[3] = 2.727"
syn_tco26 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[4] = 2.639"
syn_tco27 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[5] = 2.642"
syn_tco28 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[6] = 2.633"
syn_tco29 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[7] = 2.654"
syn_tco30 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[8] = 2.578"
syn_tco31 = " CRYPTO_HCLK->CRYPTO_AHB_M_HADDR[9] = 2.606"
syn_tco32 = " CRYPTO_HCLK->CRYPTO_AHB_M_HSIZE[0] = 2.546"
syn_tco33 = " CRYPTO_HCLK->CRYPTO_AHB_M_HSIZE[1] = 2.554"
syn_tco34 = " CRYPTO_HCLK->CRYPTO_AHB_M_HTRANS[0] = 2.818"
syn_tco35 = " CRYPTO_HCLK->CRYPTO_AHB_M_HTRANS[1] = 2.836"
syn_tco36 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[0] = 2.549"
syn_tco37 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[10] = 2.530"
syn_tco38 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[11] = 2.503"
syn_tco39 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[12] = 2.518"
syn_tco40 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[13] = 2.494"
syn_tco41 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[14] = 2.536"
syn_tco42 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[15] = 2.588"
syn_tco43 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[16] = 2.608"
syn_tco44 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[17] = 2.517"
syn_tco45 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[18] = 2.507"
syn_tco46 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[19] = 2.565"
syn_tco47 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[1] = 2.547"
syn_tco48 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[20] = 2.506"
syn_tco49 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[21] = 2.592"
syn_tco50 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[22] = 2.530"
syn_tco51 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[23] = 2.557"
syn_tco52 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[24] = 2.596"
syn_tco53 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[25] = 2.518"
syn_tco54 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[26] = 2.501"
syn_tco55 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[27] = 2.533"
syn_tco56 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[28] = 2.510"
syn_tco57 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[29] = 2.530"
syn_tco58 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[2] = 2.559"
syn_tco59 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[30] = 2.511"
syn_tco60 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[31] = 2.532"
syn_tco61 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[3] = 2.556"
syn_tco62 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[4] = 2.559"
syn_tco63 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[5] = 2.542"
syn_tco64 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[6] = 2.536"
syn_tco65 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[7] = 2.541"
syn_tco66 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[8] = 2.519"
syn_tco67 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWDATA[9] = 2.502"
syn_tco68 = " CRYPTO_HCLK->CRYPTO_AHB_M_HWRITE = 2.684"
syn_tco69 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[0] = 2.643"
syn_tco70 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[10] = 2.648"
syn_tco71 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[11] = 2.649"
syn_tco72 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[12] = 2.646"
syn_tco73 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[13] = 2.693"
syn_tco74 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[14] = 2.650"
syn_tco75 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[15] = 2.638"
syn_tco76 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[16] = 2.677"
syn_tco77 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[17] = 2.697"
syn_tco78 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[18] = 2.627"
syn_tco79 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[19] = 2.633"
syn_tco80 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[1] = 2.599"
syn_tco81 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[20] = 2.683"
syn_tco82 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[21] = 2.675"
syn_tco83 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[22] = 2.661"
syn_tco84 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[23] = 2.730"
syn_tco85 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[24] = 2.650"
syn_tco86 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[25] = 2.631"
syn_tco87 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[26] = 2.729"
syn_tco88 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[27] = 2.634"
syn_tco89 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[28] = 2.731"
syn_tco90 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[29] = 2.652"
syn_tco91 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[2] = 2.593"
syn_tco92 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[30] = 2.609"
syn_tco93 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[31] = 2.692"
syn_tco94 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[3] = 2.575"
syn_tco95 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[4] = 2.573"
syn_tco96 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[5] = 2.571"
syn_tco97 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[6] = 2.548"
syn_tco98 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[7] = 2.681"
syn_tco99 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[8] = 2.705"
syn_tco100 = " CRYPTO_HCLK->CRYPTO_AHB_S_HRDATA[9] = 2.727"
syn_tco101 = " CRYPTO_HCLK->CRYPTO_AHB_S_HREADYOUT = 2.743"
syn_tco102 = " CRYPTO_HCLK->CRYPTO_ALARM_M2F = 3.139"
syn_tco103 = " CRYPTO_HCLK->CRYPTO_BUSERROR_M2F = 2.189"
syn_tco104 = " CRYPTO_HCLK->CRYPTO_BUSY_M2F = 3.026"
syn_tco105 = " CRYPTO_HCLK->CRYPTO_COMPLETE_M2F = 3.027"
syn_tco106 = " CRYPTO_HCLK->CRYPTO_XINACCEPT_M2F = 2.510"
syn_tco107 = " CRYPTO_HCLK->CRYPTO_XRADDR_M2F[0] = 2.715"
syn_tco108 = " CRYPTO_HCLK->CRYPTO_XRADDR_M2F[1] = 2.853"
syn_tco109 = " CRYPTO_HCLK->CRYPTO_XRADDR_M2F[2] = 2.711"
syn_tco110 = " CRYPTO_HCLK->CRYPTO_XRADDR_M2F[3] = 2.667"
syn_tco111 = " CRYPTO_HCLK->CRYPTO_XRADDR_M2F[4] = 2.646"
syn_tco112 = " CRYPTO_HCLK->CRYPTO_XRADDR_M2F[5] = 2.721"
syn_tco113 = " CRYPTO_HCLK->CRYPTO_XRADDR_M2F[6] = 2.691"
syn_tco114 = " CRYPTO_HCLK->CRYPTO_XRADDR_M2F[7] = 2.692"
syn_tco115 = " CRYPTO_HCLK->CRYPTO_XRADDR_M2F[8] = 2.701"
syn_tco116 = " CRYPTO_HCLK->CRYPTO_XRADDR_M2F[9] = 2.685"
syn_tco117 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[0] = 2.579"
syn_tco118 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[10] = 2.543"
syn_tco119 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[11] = 2.559"
syn_tco120 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[12] = 2.551"
syn_tco121 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[13] = 2.539"
syn_tco122 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[14] = 2.535"
syn_tco123 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[15] = 2.473"
syn_tco124 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[16] = 2.524"
syn_tco125 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[17] = 2.467"
syn_tco126 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[18] = 2.518"
syn_tco127 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[19] = 2.520"
syn_tco128 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[1] = 2.510"
syn_tco129 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[20] = 2.502"
syn_tco130 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[21] = 2.465"
syn_tco131 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[22] = 2.460"
syn_tco132 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[23] = 2.537"
syn_tco133 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[24] = 2.541"
syn_tco134 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[25] = 2.549"
syn_tco135 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[26] = 2.523"
syn_tco136 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[27] = 2.523"
syn_tco137 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[28] = 2.524"
syn_tco138 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[29] = 2.456"
syn_tco139 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[2] = 2.529"
syn_tco140 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[30] = 2.507"
syn_tco141 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[31] = 2.521"
syn_tco142 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[3] = 2.552"
syn_tco143 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[4] = 2.491"
syn_tco144 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[5] = 2.494"
syn_tco145 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[6] = 2.514"
syn_tco146 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[7] = 2.468"
syn_tco147 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[8] = 2.453"
syn_tco148 = " CRYPTO_HCLK->CRYPTO_XRDATA_M2F[9] = 2.447"
syn_tco149 = " CRYPTO_HCLK->CRYPTO_XVALIDOUT_M2F = 2.548"
syn_tco150 = " CRYPTO_HCLK->CRYPTO_XWADDR_M2F[0] = 2.783"
syn_tco151 = " CRYPTO_HCLK->CRYPTO_XWADDR_M2F[1] = 2.774"
syn_tco152 = " CRYPTO_HCLK->CRYPTO_XWADDR_M2F[2] = 2.757"
syn_tco153 = " CRYPTO_HCLK->CRYPTO_XWADDR_M2F[3] = 2.785"
syn_tco154 = " CRYPTO_HCLK->CRYPTO_XWADDR_M2F[4] = 2.759"
syn_tco155 = " CRYPTO_HCLK->CRYPTO_XWADDR_M2F[5] = 2.718"
syn_tco156 = " CRYPTO_HCLK->CRYPTO_XWADDR_M2F[6] = 2.701"
syn_tco157 = " CRYPTO_HCLK->CRYPTO_XWADDR_M2F[7] = 2.699"
syn_tco158 = " CRYPTO_HCLK->CRYPTO_XWADDR_M2F[8] = 2.731"
syn_tco159 = " CRYPTO_HCLK->CRYPTO_XWADDR_M2F[9] = 2.739"
syn_tco160 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[0] = 0.935"
syn_tco161 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[10] = 0.973"
syn_tco162 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[11] = 0.971"
syn_tco163 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[12] = 1.040"
syn_tco164 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[13] = 1.038"
syn_tco165 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[14] = 1.037"
syn_tco166 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[15] = 1.045"
syn_tco167 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[16] = 1.037"
syn_tco168 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[17] = 1.025"
syn_tco169 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[18] = 0.968"
syn_tco170 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[19] = 1.044"
syn_tco171 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[1] = 0.942"
syn_tco172 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[20] = 1.023"
syn_tco173 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[21] = 0.939"
syn_tco174 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[22] = 1.067"
syn_tco175 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[23] = 1.031"
syn_tco176 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[24] = 0.964"
syn_tco177 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[25] = 1.013"
syn_tco178 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[26] = 1.014"
syn_tco179 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[27] = 1.014"
syn_tco180 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[28] = 0.971"
syn_tco181 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[29] = 1.035"
syn_tco182 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[2] = 0.966"
syn_tco183 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[30] = 1.062"
syn_tco184 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[31] = 0.999"
syn_tco185 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[32] = 0.949"
syn_tco186 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[33] = 0.958"
syn_tco187 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[34] = 0.994"
syn_tco188 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[35] = 1.001"
syn_tco189 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[36] = 0.988"
syn_tco190 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[37] = 1.033"
syn_tco191 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[3] = 0.960"
syn_tco192 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[4] = 0.938"
syn_tco193 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[5] = 0.992"
syn_tco194 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[6] = 0.935"
syn_tco195 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[7] = 0.996"
syn_tco196 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[8] = 1.053"
syn_tco197 = " FIC_0_ACLK->FIC_0_AXI4_M_ARADDR[9] = 1.046"
syn_tco198 = " FIC_0_ACLK->FIC_0_AXI4_M_ARBURST[0] = 1.049"
syn_tco199 = " FIC_0_ACLK->FIC_0_AXI4_M_ARBURST[1] = 0.969"
syn_tco200 = " FIC_0_ACLK->FIC_0_AXI4_M_ARCACHE[0] = 0.942"
syn_tco201 = " FIC_0_ACLK->FIC_0_AXI4_M_ARCACHE[1] = 0.950"
syn_tco202 = " FIC_0_ACLK->FIC_0_AXI4_M_ARCACHE[2] = 0.974"
syn_tco203 = " FIC_0_ACLK->FIC_0_AXI4_M_ARCACHE[3] = 0.944"
syn_tco204 = " FIC_0_ACLK->FIC_0_AXI4_M_ARID[0] = 1.021"
syn_tco205 = " FIC_0_ACLK->FIC_0_AXI4_M_ARID[1] = 1.008"
syn_tco206 = " FIC_0_ACLK->FIC_0_AXI4_M_ARID[2] = 0.952"
syn_tco207 = " FIC_0_ACLK->FIC_0_AXI4_M_ARID[3] = 1.047"
syn_tco208 = " FIC_0_ACLK->FIC_0_AXI4_M_ARID[4] = 1.035"
syn_tco209 = " FIC_0_ACLK->FIC_0_AXI4_M_ARID[5] = 0.993"
syn_tco210 = " FIC_0_ACLK->FIC_0_AXI4_M_ARID[6] = 0.972"
syn_tco211 = " FIC_0_ACLK->FIC_0_AXI4_M_ARID[7] = 0.970"
syn_tco212 = " FIC_0_ACLK->FIC_0_AXI4_M_ARLEN[0] = 1.052"
syn_tco213 = " FIC_0_ACLK->FIC_0_AXI4_M_ARLEN[1] = 1.030"
syn_tco214 = " FIC_0_ACLK->FIC_0_AXI4_M_ARLEN[2] = 1.063"
syn_tco215 = " FIC_0_ACLK->FIC_0_AXI4_M_ARLEN[3] = 1.036"
syn_tco216 = " FIC_0_ACLK->FIC_0_AXI4_M_ARLEN[4] = 0.986"
syn_tco217 = " FIC_0_ACLK->FIC_0_AXI4_M_ARLEN[5] = 0.996"
syn_tco218 = " FIC_0_ACLK->FIC_0_AXI4_M_ARLEN[6] = 1.001"
syn_tco219 = " FIC_0_ACLK->FIC_0_AXI4_M_ARLEN[7] = 1.042"
syn_tco220 = " FIC_0_ACLK->FIC_0_AXI4_M_ARLOCK = 1.022"
syn_tco221 = " FIC_0_ACLK->FIC_0_AXI4_M_ARPROT[0] = 1.009"
syn_tco222 = " FIC_0_ACLK->FIC_0_AXI4_M_ARPROT[1] = 0.944"
syn_tco223 = " FIC_0_ACLK->FIC_0_AXI4_M_ARPROT[2] = 0.955"
syn_tco224 = " FIC_0_ACLK->FIC_0_AXI4_M_ARQOS[0] = 1.031"
syn_tco225 = " FIC_0_ACLK->FIC_0_AXI4_M_ARQOS[1] = 0.971"
syn_tco226 = " FIC_0_ACLK->FIC_0_AXI4_M_ARQOS[2] = 0.969"
syn_tco227 = " FIC_0_ACLK->FIC_0_AXI4_M_ARQOS[3] = 0.895"
syn_tco228 = " FIC_0_ACLK->FIC_0_AXI4_M_ARSIZE[0] = 0.972"
syn_tco229 = " FIC_0_ACLK->FIC_0_AXI4_M_ARSIZE[1] = 1.021"
syn_tco230 = " FIC_0_ACLK->FIC_0_AXI4_M_ARSIZE[2] = 0.954"
syn_tco231 = " FIC_0_ACLK->FIC_0_AXI4_M_ARVALID = 0.790"
syn_tco232 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[0] = 0.939"
syn_tco233 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[10] = 1.006"
syn_tco234 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[11] = 1.001"
syn_tco235 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[12] = 1.000"
syn_tco236 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[13] = 0.986"
syn_tco237 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[14] = 1.003"
syn_tco238 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[15] = 0.978"
syn_tco239 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[16] = 0.960"
syn_tco240 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[17] = 1.041"
syn_tco241 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[18] = 1.010"
syn_tco242 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[19] = 0.898"
syn_tco243 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[1] = 0.915"
syn_tco244 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[20] = 1.042"
syn_tco245 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[21] = 1.041"
syn_tco246 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[22] = 0.954"
syn_tco247 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[23] = 0.985"
syn_tco248 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[24] = 1.057"
syn_tco249 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[25] = 0.985"
syn_tco250 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[26] = 0.971"
syn_tco251 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[27] = 0.946"
syn_tco252 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[28] = 1.004"
syn_tco253 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[29] = 0.936"
syn_tco254 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[2] = 0.928"
syn_tco255 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[30] = 1.023"
syn_tco256 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[31] = 1.002"
syn_tco257 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[32] = 1.016"
syn_tco258 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[33] = 1.010"
syn_tco259 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[34] = 0.906"
syn_tco260 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[35] = 0.912"
syn_tco261 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[36] = 0.976"
syn_tco262 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[37] = 0.988"
syn_tco263 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[3] = 0.923"
syn_tco264 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[4] = 0.922"
syn_tco265 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[5] = 0.888"
syn_tco266 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[6] = 0.954"
syn_tco267 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[7] = 0.966"
syn_tco268 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[8] = 0.992"
syn_tco269 = " FIC_0_ACLK->FIC_0_AXI4_M_AWADDR[9] = 0.954"
syn_tco270 = " FIC_0_ACLK->FIC_0_AXI4_M_AWBURST[0] = 0.937"
syn_tco271 = " FIC_0_ACLK->FIC_0_AXI4_M_AWBURST[1] = 0.887"
syn_tco272 = " FIC_0_ACLK->FIC_0_AXI4_M_AWCACHE[0] = 0.848"
syn_tco273 = " FIC_0_ACLK->FIC_0_AXI4_M_AWCACHE[1] = 0.921"
syn_tco274 = " FIC_0_ACLK->FIC_0_AXI4_M_AWCACHE[2] = 0.898"
syn_tco275 = " FIC_0_ACLK->FIC_0_AXI4_M_AWCACHE[3] = 0.899"
syn_tco276 = " FIC_0_ACLK->FIC_0_AXI4_M_AWID[0] = 0.948"
syn_tco277 = " FIC_0_ACLK->FIC_0_AXI4_M_AWID[1] = 0.948"
syn_tco278 = " FIC_0_ACLK->FIC_0_AXI4_M_AWID[2] = 0.943"
syn_tco279 = " FIC_0_ACLK->FIC_0_AXI4_M_AWID[3] = 0.954"
syn_tco280 = " FIC_0_ACLK->FIC_0_AXI4_M_AWID[4] = 0.930"
syn_tco281 = " FIC_0_ACLK->FIC_0_AXI4_M_AWID[5] = 0.945"
syn_tco282 = " FIC_0_ACLK->FIC_0_AXI4_M_AWID[6] = 0.915"
syn_tco283 = " FIC_0_ACLK->FIC_0_AXI4_M_AWID[7] = 0.885"
syn_tco284 = " FIC_0_ACLK->FIC_0_AXI4_M_AWLEN[0] = 0.833"
syn_tco285 = " FIC_0_ACLK->FIC_0_AXI4_M_AWLEN[1] = 0.823"
syn_tco286 = " FIC_0_ACLK->FIC_0_AXI4_M_AWLEN[2] = 0.887"
syn_tco287 = " FIC_0_ACLK->FIC_0_AXI4_M_AWLEN[3] = 0.854"
syn_tco288 = " FIC_0_ACLK->FIC_0_AXI4_M_AWLEN[4] = 0.861"
syn_tco289 = " FIC_0_ACLK->FIC_0_AXI4_M_AWLEN[5] = 0.895"
syn_tco290 = " FIC_0_ACLK->FIC_0_AXI4_M_AWLEN[6] = 0.903"
syn_tco291 = " FIC_0_ACLK->FIC_0_AXI4_M_AWLEN[7] = 0.888"
syn_tco292 = " FIC_0_ACLK->FIC_0_AXI4_M_AWLOCK = 0.828"
syn_tco293 = " FIC_0_ACLK->FIC_0_AXI4_M_AWPROT[0] = 0.881"
syn_tco294 = " FIC_0_ACLK->FIC_0_AXI4_M_AWPROT[1] = 0.883"
syn_tco295 = " FIC_0_ACLK->FIC_0_AXI4_M_AWPROT[2] = 0.844"
syn_tco296 = " FIC_0_ACLK->FIC_0_AXI4_M_AWQOS[0] = 0.848"
syn_tco297 = " FIC_0_ACLK->FIC_0_AXI4_M_AWQOS[1] = 0.919"
syn_tco298 = " FIC_0_ACLK->FIC_0_AXI4_M_AWQOS[2] = 0.859"
syn_tco299 = " FIC_0_ACLK->FIC_0_AXI4_M_AWQOS[3] = 0.863"
syn_tco300 = " FIC_0_ACLK->FIC_0_AXI4_M_AWSIZE[0] = 0.850"
syn_tco301 = " FIC_0_ACLK->FIC_0_AXI4_M_AWSIZE[1] = 0.895"
syn_tco302 = " FIC_0_ACLK->FIC_0_AXI4_M_AWSIZE[2] = 0.814"
syn_tco303 = " FIC_0_ACLK->FIC_0_AXI4_M_AWVALID = 0.534"
syn_tco304 = " FIC_0_ACLK->FIC_0_AXI4_M_BREADY = 0.651"
syn_tco305 = " FIC_0_ACLK->FIC_0_AXI4_M_RREADY = 0.596"
syn_tco306 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[0] = 0.900"
syn_tco307 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[10] = 0.891"
syn_tco308 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[11] = 0.884"
syn_tco309 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[12] = 0.937"
syn_tco310 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[13] = 0.880"
syn_tco311 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[14] = 0.885"
syn_tco312 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[15] = 0.924"
syn_tco313 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[16] = 0.922"
syn_tco314 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[17] = 0.892"
syn_tco315 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[18] = 0.926"
syn_tco316 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[19] = 0.888"
syn_tco317 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[1] = 0.891"
syn_tco318 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[20] = 0.919"
syn_tco319 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[21] = 0.923"
syn_tco320 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[22] = 0.886"
syn_tco321 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[23] = 0.917"
syn_tco322 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[24] = 0.899"
syn_tco323 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[25] = 0.913"
syn_tco324 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[26] = 0.880"
syn_tco325 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[27] = 0.894"
syn_tco326 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[28] = 0.891"
syn_tco327 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[29] = 0.904"
syn_tco328 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[2] = 0.875"
syn_tco329 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[30] = 0.881"
syn_tco330 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[31] = 0.927"
syn_tco331 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[32] = 0.909"
syn_tco332 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[33] = 0.912"
syn_tco333 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[34] = 0.916"
syn_tco334 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[35] = 0.931"
syn_tco335 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[36] = 0.897"
syn_tco336 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[37] = 0.897"
syn_tco337 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[38] = 0.898"
syn_tco338 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[39] = 0.914"
syn_tco339 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[3] = 0.896"
syn_tco340 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[40] = 0.910"
syn_tco341 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[41] = 0.904"
syn_tco342 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[42] = 0.883"
syn_tco343 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[43] = 0.905"
syn_tco344 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[44] = 0.909"
syn_tco345 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[45] = 0.893"
syn_tco346 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[46] = 0.936"
syn_tco347 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[47] = 0.922"
syn_tco348 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[48] = 0.956"
syn_tco349 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[49] = 0.898"
syn_tco350 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[4] = 0.890"
syn_tco351 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[50] = 0.916"
syn_tco352 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[51] = 0.921"
syn_tco353 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[52] = 0.914"
syn_tco354 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[53] = 0.895"
syn_tco355 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[54] = 0.879"
syn_tco356 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[55] = 0.900"
syn_tco357 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[56] = 0.910"
syn_tco358 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[57] = 0.899"
syn_tco359 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[58] = 0.896"
syn_tco360 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[59] = 0.931"
syn_tco361 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[5] = 0.890"
syn_tco362 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[60] = 0.924"
syn_tco363 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[61] = 0.915"
syn_tco364 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[62] = 0.936"
syn_tco365 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[63] = 0.881"
syn_tco366 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[6] = 0.906"
syn_tco367 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[7] = 0.886"
syn_tco368 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[8] = 0.891"
syn_tco369 = " FIC_0_ACLK->FIC_0_AXI4_M_WDATA[9] = 0.901"
syn_tco370 = " FIC_0_ACLK->FIC_0_AXI4_M_WLAST = 0.891"
syn_tco371 = " FIC_0_ACLK->FIC_0_AXI4_M_WSTRB[0] = 0.910"
syn_tco372 = " FIC_0_ACLK->FIC_0_AXI4_M_WSTRB[1] = 0.886"
syn_tco373 = " FIC_0_ACLK->FIC_0_AXI4_M_WSTRB[2] = 0.958"
syn_tco374 = " FIC_0_ACLK->FIC_0_AXI4_M_WSTRB[3] = 0.905"
syn_tco375 = " FIC_0_ACLK->FIC_0_AXI4_M_WSTRB[4] = 0.917"
syn_tco376 = " FIC_0_ACLK->FIC_0_AXI4_M_WSTRB[5] = 0.895"
syn_tco377 = " FIC_0_ACLK->FIC_0_AXI4_M_WSTRB[6] = 0.933"
syn_tco378 = " FIC_0_ACLK->FIC_0_AXI4_M_WSTRB[7] = 0.886"
syn_tco379 = " FIC_0_ACLK->FIC_0_AXI4_M_WVALID = 0.572"
syn_tco380 = " FIC_0_ACLK->FIC_0_AXI4_S_ARREADY = 0.913"
syn_tco381 = " FIC_0_ACLK->FIC_0_AXI4_S_AWREADY = 0.832"
syn_tco382 = " FIC_0_ACLK->FIC_0_AXI4_S_BID[0] = 1.035"
syn_tco383 = " FIC_0_ACLK->FIC_0_AXI4_S_BID[1] = 1.024"
syn_tco384 = " FIC_0_ACLK->FIC_0_AXI4_S_BID[2] = 1.033"
syn_tco385 = " FIC_0_ACLK->FIC_0_AXI4_S_BID[3] = 1.005"
syn_tco386 = " FIC_0_ACLK->FIC_0_AXI4_S_BRESP[0] = 1.023"
syn_tco387 = " FIC_0_ACLK->FIC_0_AXI4_S_BRESP[1] = 0.956"
syn_tco388 = " FIC_0_ACLK->FIC_0_AXI4_S_BVALID = 0.803"
syn_tco389 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[0] = 0.917"
syn_tco390 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[10] = 0.953"
syn_tco391 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[11] = 0.953"
syn_tco392 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[12] = 0.971"
syn_tco393 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[13] = 0.981"
syn_tco394 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[14] = 0.996"
syn_tco395 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[15] = 0.920"
syn_tco396 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[16] = 1.000"
syn_tco397 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[17] = 0.943"
syn_tco398 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[18] = 0.927"
syn_tco399 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[19] = 0.934"
syn_tco400 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[1] = 0.950"
syn_tco401 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[20] = 0.978"
syn_tco402 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[21] = 1.011"
syn_tco403 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[22] = 0.929"
syn_tco404 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[23] = 0.896"
syn_tco405 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[24] = 0.958"
syn_tco406 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[25] = 0.954"
syn_tco407 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[26] = 0.895"
syn_tco408 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[27] = 0.930"
syn_tco409 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[28] = 0.940"
syn_tco410 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[29] = 0.912"
syn_tco411 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[2] = 1.023"
syn_tco412 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[30] = 0.923"
syn_tco413 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[31] = 0.934"
syn_tco414 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[32] = 0.928"
syn_tco415 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[33] = 0.962"
syn_tco416 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[34] = 0.939"
syn_tco417 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[35] = 0.934"
syn_tco418 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[36] = 0.969"
syn_tco419 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[37] = 0.916"
syn_tco420 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[38] = 0.980"
syn_tco421 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[39] = 0.947"
syn_tco422 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[3] = 0.984"
syn_tco423 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[40] = 0.972"
syn_tco424 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[41] = 0.977"
syn_tco425 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[42] = 1.015"
syn_tco426 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[43] = 0.936"
syn_tco427 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[44] = 0.957"
syn_tco428 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[45] = 0.967"
syn_tco429 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[46] = 0.926"
syn_tco430 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[47] = 0.953"
syn_tco431 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[48] = 0.964"
syn_tco432 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[49] = 0.973"
syn_tco433 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[4] = 0.967"
syn_tco434 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[50] = 0.983"
syn_tco435 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[51] = 0.914"
syn_tco436 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[52] = 0.948"
syn_tco437 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[53] = 0.908"
syn_tco438 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[54] = 0.928"
syn_tco439 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[55] = 0.926"
syn_tco440 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[56] = 0.971"
syn_tco441 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[57] = 0.968"
syn_tco442 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[58] = 0.890"
syn_tco443 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[59] = 0.944"
syn_tco444 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[5] = 0.953"
syn_tco445 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[60] = 0.966"
syn_tco446 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[61] = 0.921"
syn_tco447 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[62] = 0.887"
syn_tco448 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[63] = 1.021"
syn_tco449 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[6] = 1.026"
syn_tco450 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[7] = 0.976"
syn_tco451 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[8] = 0.974"
syn_tco452 = " FIC_0_ACLK->FIC_0_AXI4_S_RDATA[9] = 0.979"
syn_tco453 = " FIC_0_ACLK->FIC_0_AXI4_S_RID[0] = 0.945"
syn_tco454 = " FIC_0_ACLK->FIC_0_AXI4_S_RID[1] = 0.981"
syn_tco455 = " FIC_0_ACLK->FIC_0_AXI4_S_RID[2] = 0.990"
syn_tco456 = " FIC_0_ACLK->FIC_0_AXI4_S_RID[3] = 0.982"
syn_tco457 = " FIC_0_ACLK->FIC_0_AXI4_S_RLAST = 1.009"
syn_tco458 = " FIC_0_ACLK->FIC_0_AXI4_S_RRESP[0] = 0.987"
syn_tco459 = " FIC_0_ACLK->FIC_0_AXI4_S_RRESP[1] = 0.966"
syn_tco460 = " FIC_0_ACLK->FIC_0_AXI4_S_RVALID = 0.868"
syn_tco461 = " FIC_0_ACLK->FIC_0_AXI4_S_WREADY = 0.859"
syn_tco462 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[0] = 0.969"
syn_tco463 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[10] = 0.967"
syn_tco464 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[11] = 0.980"
syn_tco465 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[12] = 0.925"
syn_tco466 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[13] = 0.933"
syn_tco467 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[14] = 0.963"
syn_tco468 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[15] = 0.963"
syn_tco469 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[16] = 0.949"
syn_tco470 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[17] = 0.940"
syn_tco471 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[18] = 0.980"
syn_tco472 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[19] = 0.982"
syn_tco473 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[1] = 0.939"
syn_tco474 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[20] = 1.005"
syn_tco475 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[21] = 0.998"
syn_tco476 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[22] = 0.996"
syn_tco477 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[23] = 0.990"
syn_tco478 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[24] = 0.994"
syn_tco479 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[25] = 1.016"
syn_tco480 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[26] = 1.001"
syn_tco481 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[27] = 0.977"
syn_tco482 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[28] = 0.973"
syn_tco483 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[29] = 0.973"
syn_tco484 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[2] = 0.974"
syn_tco485 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[30] = 0.969"
syn_tco486 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[31] = 0.971"
syn_tco487 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[32] = 1.006"
syn_tco488 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[33] = 1.036"
syn_tco489 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[34] = 1.014"
syn_tco490 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[35] = 0.942"
syn_tco491 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[36] = 0.979"
syn_tco492 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[37] = 0.907"
syn_tco493 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[3] = 0.950"
syn_tco494 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[4] = 0.938"
syn_tco495 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[5] = 0.960"
syn_tco496 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[6] = 0.980"
syn_tco497 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[7] = 0.990"
syn_tco498 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[8] = 0.969"
syn_tco499 = " FIC_1_ACLK->FIC_1_AXI4_M_ARADDR[9] = 0.990"
syn_tco500 = " FIC_1_ACLK->FIC_1_AXI4_M_ARBURST[0] = 0.977"
syn_tco501 = " FIC_1_ACLK->FIC_1_AXI4_M_ARBURST[1] = 0.982"
syn_tco502 = " FIC_1_ACLK->FIC_1_AXI4_M_ARCACHE[0] = 0.944"
syn_tco503 = " FIC_1_ACLK->FIC_1_AXI4_M_ARCACHE[1] = 0.899"
syn_tco504 = " FIC_1_ACLK->FIC_1_AXI4_M_ARCACHE[2] = 0.850"
syn_tco505 = " FIC_1_ACLK->FIC_1_AXI4_M_ARCACHE[3] = 0.845"
syn_tco506 = " FIC_1_ACLK->FIC_1_AXI4_M_ARID[0] = 0.909"
syn_tco507 = " FIC_1_ACLK->FIC_1_AXI4_M_ARID[1] = 0.950"
syn_tco508 = " FIC_1_ACLK->FIC_1_AXI4_M_ARID[2] = 0.925"
syn_tco509 = " FIC_1_ACLK->FIC_1_AXI4_M_ARID[3] = 1.018"
syn_tco510 = " FIC_1_ACLK->FIC_1_AXI4_M_ARID[4] = 0.975"
syn_tco511 = " FIC_1_ACLK->FIC_1_AXI4_M_ARID[5] = 0.964"
syn_tco512 = " FIC_1_ACLK->FIC_1_AXI4_M_ARID[6] = 0.973"
syn_tco513 = " FIC_1_ACLK->FIC_1_AXI4_M_ARID[7] = 0.986"
syn_tco514 = " FIC_1_ACLK->FIC_1_AXI4_M_ARLEN[0] = 0.889"
syn_tco515 = " FIC_1_ACLK->FIC_1_AXI4_M_ARLEN[1] = 0.979"
syn_tco516 = " FIC_1_ACLK->FIC_1_AXI4_M_ARLEN[2] = 0.962"
syn_tco517 = " FIC_1_ACLK->FIC_1_AXI4_M_ARLEN[3] = 0.965"
syn_tco518 = " FIC_1_ACLK->FIC_1_AXI4_M_ARLEN[4] = 0.988"
syn_tco519 = " FIC_1_ACLK->FIC_1_AXI4_M_ARLEN[5] = 0.990"
syn_tco520 = " FIC_1_ACLK->FIC_1_AXI4_M_ARLEN[6] = 0.980"
syn_tco521 = " FIC_1_ACLK->FIC_1_AXI4_M_ARLEN[7] = 0.965"
syn_tco522 = " FIC_1_ACLK->FIC_1_AXI4_M_ARLOCK = 0.971"
syn_tco523 = " FIC_1_ACLK->FIC_1_AXI4_M_ARPROT[0] = 1.010"
syn_tco524 = " FIC_1_ACLK->FIC_1_AXI4_M_ARPROT[1] = 0.977"
syn_tco525 = " FIC_1_ACLK->FIC_1_AXI4_M_ARPROT[2] = 0.978"
syn_tco526 = " FIC_1_ACLK->FIC_1_AXI4_M_ARQOS[0] = 1.013"
syn_tco527 = " FIC_1_ACLK->FIC_1_AXI4_M_ARQOS[1] = 0.963"
syn_tco528 = " FIC_1_ACLK->FIC_1_AXI4_M_ARQOS[2] = 0.999"
syn_tco529 = " FIC_1_ACLK->FIC_1_AXI4_M_ARQOS[3] = 0.972"
syn_tco530 = " FIC_1_ACLK->FIC_1_AXI4_M_ARSIZE[0] = 0.993"
syn_tco531 = " FIC_1_ACLK->FIC_1_AXI4_M_ARSIZE[1] = 0.993"
syn_tco532 = " FIC_1_ACLK->FIC_1_AXI4_M_ARSIZE[2] = 0.997"
syn_tco533 = " FIC_1_ACLK->FIC_1_AXI4_M_ARVALID = 0.670"
syn_tco534 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[0] = 0.812"
syn_tco535 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[10] = 0.858"
syn_tco536 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[11] = 0.796"
syn_tco537 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[12] = 0.797"
syn_tco538 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[13] = 0.781"
syn_tco539 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[14] = 0.786"
syn_tco540 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[15] = 0.833"
syn_tco541 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[16] = 0.831"
syn_tco542 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[17] = 0.884"
syn_tco543 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[18] = 0.884"
syn_tco544 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[19] = 0.921"
syn_tco545 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[1] = 0.895"
syn_tco546 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[20] = 0.922"
syn_tco547 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[21] = 0.924"
syn_tco548 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[22] = 0.924"
syn_tco549 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[23] = 0.838"
syn_tco550 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[24] = 0.939"
syn_tco551 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[25] = 0.874"
syn_tco552 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[26] = 0.887"
syn_tco553 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[27] = 0.869"
syn_tco554 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[28] = 0.892"
syn_tco555 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[29] = 0.886"
syn_tco556 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[2] = 0.837"
syn_tco557 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[30] = 0.906"
syn_tco558 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[31] = 0.826"
syn_tco559 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[32] = 0.838"
syn_tco560 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[33] = 0.845"
syn_tco561 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[34] = 0.808"
syn_tco562 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[35] = 0.822"
syn_tco563 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[36] = 0.844"
syn_tco564 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[37] = 0.876"
syn_tco565 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[3] = 0.860"
syn_tco566 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[4] = 0.874"
syn_tco567 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[5] = 0.850"
syn_tco568 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[6] = 0.840"
syn_tco569 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[7] = 0.866"
syn_tco570 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[8] = 0.849"
syn_tco571 = " FIC_1_ACLK->FIC_1_AXI4_M_AWADDR[9] = 0.880"
syn_tco572 = " FIC_1_ACLK->FIC_1_AXI4_M_AWBURST[0] = 0.849"
syn_tco573 = " FIC_1_ACLK->FIC_1_AXI4_M_AWBURST[1] = 0.839"
syn_tco574 = " FIC_1_ACLK->FIC_1_AXI4_M_AWCACHE[0] = 0.835"
syn_tco575 = " FIC_1_ACLK->FIC_1_AXI4_M_AWCACHE[1] = 0.864"
syn_tco576 = " FIC_1_ACLK->FIC_1_AXI4_M_AWCACHE[2] = 0.853"
syn_tco577 = " FIC_1_ACLK->FIC_1_AXI4_M_AWCACHE[3] = 0.846"
syn_tco578 = " FIC_1_ACLK->FIC_1_AXI4_M_AWID[0] = 0.857"
syn_tco579 = " FIC_1_ACLK->FIC_1_AXI4_M_AWID[1] = 0.715"
syn_tco580 = " FIC_1_ACLK->FIC_1_AXI4_M_AWID[2] = 0.704"
syn_tco581 = " FIC_1_ACLK->FIC_1_AXI4_M_AWID[3] = 0.708"
syn_tco582 = " FIC_1_ACLK->FIC_1_AXI4_M_AWID[4] = 0.841"
syn_tco583 = " FIC_1_ACLK->FIC_1_AXI4_M_AWID[5] = 0.761"
syn_tco584 = " FIC_1_ACLK->FIC_1_AXI4_M_AWID[6] = 0.766"
syn_tco585 = " FIC_1_ACLK->FIC_1_AXI4_M_AWID[7] = 0.728"
syn_tco586 = " FIC_1_ACLK->FIC_1_AXI4_M_AWLEN[0] = 0.849"
syn_tco587 = " FIC_1_ACLK->FIC_1_AXI4_M_AWLEN[1] = 0.865"
syn_tco588 = " FIC_1_ACLK->FIC_1_AXI4_M_AWLEN[2] = 0.875"
syn_tco589 = " FIC_1_ACLK->FIC_1_AXI4_M_AWLEN[3] = 0.840"
syn_tco590 = " FIC_1_ACLK->FIC_1_AXI4_M_AWLEN[4] = 0.873"
syn_tco591 = " FIC_1_ACLK->FIC_1_AXI4_M_AWLEN[5] = 0.855"
syn_tco592 = " FIC_1_ACLK->FIC_1_AXI4_M_AWLEN[6] = 0.845"
syn_tco593 = " FIC_1_ACLK->FIC_1_AXI4_M_AWLEN[7] = 0.819"
syn_tco594 = " FIC_1_ACLK->FIC_1_AXI4_M_AWLOCK = 0.848"
syn_tco595 = " FIC_1_ACLK->FIC_1_AXI4_M_AWPROT[0] = 0.876"
syn_tco596 = " FIC_1_ACLK->FIC_1_AXI4_M_AWPROT[1] = 0.863"
syn_tco597 = " FIC_1_ACLK->FIC_1_AXI4_M_AWPROT[2] = 0.850"
syn_tco598 = " FIC_1_ACLK->FIC_1_AXI4_M_AWQOS[0] = 0.810"
syn_tco599 = " FIC_1_ACLK->FIC_1_AXI4_M_AWQOS[1] = 0.849"
syn_tco600 = " FIC_1_ACLK->FIC_1_AXI4_M_AWQOS[2] = 0.835"
syn_tco601 = " FIC_1_ACLK->FIC_1_AXI4_M_AWQOS[3] = 0.853"
syn_tco602 = " FIC_1_ACLK->FIC_1_AXI4_M_AWSIZE[0] = 0.842"
syn_tco603 = " FIC_1_ACLK->FIC_1_AXI4_M_AWSIZE[1] = 0.883"
syn_tco604 = " FIC_1_ACLK->FIC_1_AXI4_M_AWSIZE[2] = 0.880"
syn_tco605 = " FIC_1_ACLK->FIC_1_AXI4_M_AWVALID = 0.398"
syn_tco606 = " FIC_1_ACLK->FIC_1_AXI4_M_BREADY = 0.630"
syn_tco607 = " FIC_1_ACLK->FIC_1_AXI4_M_RREADY = 0.609"
syn_tco608 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[0] = 0.913"
syn_tco609 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[10] = 0.912"
syn_tco610 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[11] = 0.894"
syn_tco611 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[12] = 0.895"
syn_tco612 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[13] = 0.878"
syn_tco613 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[14] = 0.896"
syn_tco614 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[15] = 0.898"
syn_tco615 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[16] = 0.905"
syn_tco616 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[17] = 0.903"
syn_tco617 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[18] = 0.898"
syn_tco618 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[19] = 0.899"
syn_tco619 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[1] = 0.909"
syn_tco620 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[20] = 0.895"
syn_tco621 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[21] = 0.898"
syn_tco622 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[22] = 0.879"
syn_tco623 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[23] = 0.885"
syn_tco624 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[24] = 0.861"
syn_tco625 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[25] = 0.870"
syn_tco626 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[26] = 0.884"
syn_tco627 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[27] = 0.861"
syn_tco628 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[28] = 0.862"
syn_tco629 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[29] = 0.929"
syn_tco630 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[2] = 0.889"
syn_tco631 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[30] = 0.852"
syn_tco632 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[31] = 0.895"
syn_tco633 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[32] = 0.895"
syn_tco634 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[33] = 0.908"
syn_tco635 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[34] = 0.925"
syn_tco636 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[35] = 0.908"
syn_tco637 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[36] = 0.908"
syn_tco638 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[37] = 0.897"
syn_tco639 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[38] = 0.923"
syn_tco640 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[39] = 0.884"
syn_tco641 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[3] = 0.926"
syn_tco642 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[40] = 0.906"
syn_tco643 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[41] = 0.949"
syn_tco644 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[42] = 0.949"
syn_tco645 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[43] = 0.886"
syn_tco646 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[44] = 0.926"
syn_tco647 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[45] = 0.889"
syn_tco648 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[46] = 0.899"
syn_tco649 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[47] = 0.909"
syn_tco650 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[48] = 0.876"
syn_tco651 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[49] = 0.884"
syn_tco652 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[4] = 0.886"
syn_tco653 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[50] = 0.869"
syn_tco654 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[51] = 0.943"
syn_tco655 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[52] = 0.953"
syn_tco656 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[53] = 0.964"
syn_tco657 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[54] = 0.956"
syn_tco658 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[55] = 0.918"
syn_tco659 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[56] = 0.910"
syn_tco660 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[57] = 0.930"
syn_tco661 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[58] = 0.933"
syn_tco662 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[59] = 0.887"
syn_tco663 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[5] = 0.886"
syn_tco664 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[60] = 0.879"
syn_tco665 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[61] = 0.874"
syn_tco666 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[62] = 0.896"
syn_tco667 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[63] = 0.855"
syn_tco668 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[6] = 0.897"
syn_tco669 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[7] = 0.882"
syn_tco670 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[8] = 0.870"
syn_tco671 = " FIC_1_ACLK->FIC_1_AXI4_M_WDATA[9] = 0.894"
syn_tco672 = " FIC_1_ACLK->FIC_1_AXI4_M_WLAST = 0.914"
syn_tco673 = " FIC_1_ACLK->FIC_1_AXI4_M_WSTRB[0] = 0.888"
syn_tco674 = " FIC_1_ACLK->FIC_1_AXI4_M_WSTRB[1] = 0.923"
syn_tco675 = " FIC_1_ACLK->FIC_1_AXI4_M_WSTRB[2] = 0.927"
syn_tco676 = " FIC_1_ACLK->FIC_1_AXI4_M_WSTRB[3] = 0.920"
syn_tco677 = " FIC_1_ACLK->FIC_1_AXI4_M_WSTRB[4] = 0.920"
syn_tco678 = " FIC_1_ACLK->FIC_1_AXI4_M_WSTRB[5] = 0.896"
syn_tco679 = " FIC_1_ACLK->FIC_1_AXI4_M_WSTRB[6] = 0.931"
syn_tco680 = " FIC_1_ACLK->FIC_1_AXI4_M_WSTRB[7] = 0.899"
syn_tco681 = " FIC_1_ACLK->FIC_1_AXI4_M_WVALID = 0.509"
syn_tco682 = " FIC_1_ACLK->FIC_1_AXI4_S_ARREADY = 0.916"
syn_tco683 = " FIC_1_ACLK->FIC_1_AXI4_S_AWREADY = 0.899"
syn_tco684 = " FIC_1_ACLK->FIC_1_AXI4_S_BID[0] = 1.007"
syn_tco685 = " FIC_1_ACLK->FIC_1_AXI4_S_BID[1] = 0.873"
syn_tco686 = " FIC_1_ACLK->FIC_1_AXI4_S_BID[2] = 0.973"
syn_tco687 = " FIC_1_ACLK->FIC_1_AXI4_S_BID[3] = 0.964"
syn_tco688 = " FIC_1_ACLK->FIC_1_AXI4_S_BRESP[0] = 0.971"
syn_tco689 = " FIC_1_ACLK->FIC_1_AXI4_S_BRESP[1] = 0.822"
syn_tco690 = " FIC_1_ACLK->FIC_1_AXI4_S_BVALID = 0.796"
syn_tco691 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[0] = 0.992"
syn_tco692 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[10] = 0.950"
syn_tco693 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[11] = 0.950"
syn_tco694 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[12] = 0.948"
syn_tco695 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[13] = 0.953"
syn_tco696 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[14] = 0.963"
syn_tco697 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[15] = 0.951"
syn_tco698 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[16] = 0.951"
syn_tco699 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[17] = 0.892"
syn_tco700 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[18] = 0.997"
syn_tco701 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[19] = 0.972"
syn_tco702 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[1] = 0.888"
syn_tco703 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[20] = 0.981"
syn_tco704 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[21] = 0.964"
syn_tco705 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[22] = 0.973"
syn_tco706 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[23] = 0.986"
syn_tco707 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[24] = 0.979"
syn_tco708 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[25] = 0.986"
syn_tco709 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[26] = 0.989"
syn_tco710 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[27] = 0.969"
syn_tco711 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[28] = 1.025"
syn_tco712 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[29] = 0.990"
syn_tco713 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[2] = 0.936"
syn_tco714 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[30] = 0.988"
syn_tco715 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[31] = 0.937"
syn_tco716 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[32] = 0.929"
syn_tco717 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[33] = 1.002"
syn_tco718 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[34] = 1.003"
syn_tco719 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[35] = 0.974"
syn_tco720 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[36] = 1.008"
syn_tco721 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[37] = 0.931"
syn_tco722 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[38] = 1.030"
syn_tco723 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[39] = 0.966"
syn_tco724 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[3] = 0.923"
syn_tco725 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[40] = 0.919"
syn_tco726 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[41] = 0.990"
syn_tco727 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[42] = 0.996"
syn_tco728 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[43] = 1.033"
syn_tco729 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[44] = 1.029"
syn_tco730 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[45] = 0.937"
syn_tco731 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[46] = 0.968"
syn_tco732 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[47] = 0.972"
syn_tco733 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[48] = 0.992"
syn_tco734 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[49] = 0.982"
syn_tco735 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[4] = 0.971"
syn_tco736 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[50] = 0.999"
syn_tco737 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[51] = 0.992"
syn_tco738 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[52] = 0.970"
syn_tco739 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[53] = 0.960"
syn_tco740 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[54] = 0.970"
syn_tco741 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[55] = 0.979"
syn_tco742 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[56] = 1.016"
syn_tco743 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[57] = 0.973"
syn_tco744 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[58] = 0.969"
syn_tco745 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[59] = 0.993"
syn_tco746 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[5] = 0.924"
syn_tco747 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[60] = 1.006"
syn_tco748 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[61] = 0.987"
syn_tco749 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[62] = 0.912"
syn_tco750 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[63] = 0.938"
syn_tco751 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[6] = 0.967"
syn_tco752 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[7] = 0.977"
syn_tco753 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[8] = 0.955"
syn_tco754 = " FIC_1_ACLK->FIC_1_AXI4_S_RDATA[9] = 0.950"
syn_tco755 = " FIC_1_ACLK->FIC_1_AXI4_S_RID[0] = 0.919"
syn_tco756 = " FIC_1_ACLK->FIC_1_AXI4_S_RID[1] = 0.953"
syn_tco757 = " FIC_1_ACLK->FIC_1_AXI4_S_RID[2] = 0.915"
syn_tco758 = " FIC_1_ACLK->FIC_1_AXI4_S_RID[3] = 0.979"
syn_tco759 = " FIC_1_ACLK->FIC_1_AXI4_S_RLAST = 0.941"
syn_tco760 = " FIC_1_ACLK->FIC_1_AXI4_S_RRESP[0] = 0.962"
syn_tco761 = " FIC_1_ACLK->FIC_1_AXI4_S_RRESP[1] = 0.949"
syn_tco762 = " FIC_1_ACLK->FIC_1_AXI4_S_RVALID = 0.573"
syn_tco763 = " FIC_1_ACLK->FIC_1_AXI4_S_WREADY = 0.766"
syn_tco764 = " FIC_2_ACLK->FIC_2_AXI4_S_ARREADY = 0.844"
syn_tco765 = " FIC_2_ACLK->FIC_2_AXI4_S_AWREADY = 0.868"
syn_tco766 = " FIC_2_ACLK->FIC_2_AXI4_S_BID[0] = 0.864"
syn_tco767 = " FIC_2_ACLK->FIC_2_AXI4_S_BID[1] = 0.857"
syn_tco768 = " FIC_2_ACLK->FIC_2_AXI4_S_BID[2] = 0.965"
syn_tco769 = " FIC_2_ACLK->FIC_2_AXI4_S_BID[3] = 0.870"
syn_tco770 = " FIC_2_ACLK->FIC_2_AXI4_S_BRESP[0] = 0.860"
syn_tco771 = " FIC_2_ACLK->FIC_2_AXI4_S_BRESP[1] = 0.892"
syn_tco772 = " FIC_2_ACLK->FIC_2_AXI4_S_BVALID = 0.718"
syn_tco773 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[0] = 0.838"
syn_tco774 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[10] = 0.831"
syn_tco775 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[11] = 0.815"
syn_tco776 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[12] = 0.812"
syn_tco777 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[13] = 0.831"
syn_tco778 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[14] = 0.841"
syn_tco779 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[15] = 0.845"
syn_tco780 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[16] = 0.847"
syn_tco781 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[17] = 0.874"
syn_tco782 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[18] = 0.947"
syn_tco783 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[19] = 0.842"
syn_tco784 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[1] = 0.832"
syn_tco785 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[20] = 0.901"
syn_tco786 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[21] = 0.835"
syn_tco787 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[22] = 0.870"
syn_tco788 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[23] = 0.879"
syn_tco789 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[24] = 0.841"
syn_tco790 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[25] = 0.879"
syn_tco791 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[26] = 0.846"
syn_tco792 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[27] = 0.925"
syn_tco793 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[28] = 0.894"
syn_tco794 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[29] = 0.844"
syn_tco795 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[2] = 0.844"
syn_tco796 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[30] = 0.892"
syn_tco797 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[31] = 0.861"
syn_tco798 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[32] = 0.878"
syn_tco799 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[33] = 0.871"
syn_tco800 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[34] = 0.865"
syn_tco801 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[35] = 0.885"
syn_tco802 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[36] = 0.868"
syn_tco803 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[37] = 0.868"
syn_tco804 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[38] = 0.857"
syn_tco805 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[39] = 0.850"
syn_tco806 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[3] = 0.858"
syn_tco807 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[40] = 0.860"
syn_tco808 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[41] = 0.867"
syn_tco809 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[42] = 0.863"
syn_tco810 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[43] = 0.905"
syn_tco811 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[44] = 0.880"
syn_tco812 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[45] = 0.889"
syn_tco813 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[46] = 0.894"
syn_tco814 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[47] = 0.889"
syn_tco815 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[48] = 0.892"
syn_tco816 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[49] = 0.882"
syn_tco817 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[4] = 0.855"
syn_tco818 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[50] = 0.879"
syn_tco819 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[51] = 0.892"
syn_tco820 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[52] = 0.893"
syn_tco821 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[53] = 0.863"
syn_tco822 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[54] = 0.875"
syn_tco823 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[55] = 0.914"
syn_tco824 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[56] = 0.948"
syn_tco825 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[57] = 0.896"
syn_tco826 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[58] = 0.887"
syn_tco827 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[59] = 0.886"
syn_tco828 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[5] = 0.825"
syn_tco829 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[60] = 0.916"
syn_tco830 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[61] = 0.853"
syn_tco831 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[62] = 0.915"
syn_tco832 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[63] = 0.893"
syn_tco833 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[6] = 0.826"
syn_tco834 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[7] = 0.835"
syn_tco835 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[8] = 0.841"
syn_tco836 = " FIC_2_ACLK->FIC_2_AXI4_S_RDATA[9] = 0.886"
syn_tco837 = " FIC_2_ACLK->FIC_2_AXI4_S_RID[0] = 0.866"
syn_tco838 = " FIC_2_ACLK->FIC_2_AXI4_S_RID[1] = 0.859"
syn_tco839 = " FIC_2_ACLK->FIC_2_AXI4_S_RID[2] = 0.811"
syn_tco840 = " FIC_2_ACLK->FIC_2_AXI4_S_RID[3] = 0.838"
syn_tco841 = " FIC_2_ACLK->FIC_2_AXI4_S_RLAST = 0.809"
syn_tco842 = " FIC_2_ACLK->FIC_2_AXI4_S_RRESP[0] = 0.842"
syn_tco843 = " FIC_2_ACLK->FIC_2_AXI4_S_RRESP[1] = 0.845"
syn_tco844 = " FIC_2_ACLK->FIC_2_AXI4_S_RVALID = 0.391"
syn_tco845 = " FIC_2_ACLK->FIC_2_AXI4_S_WREADY = 0.759"
syn_tco846 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[10] = 1.772"
syn_tco847 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[11] = 1.768"
syn_tco848 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[12] = 1.758"
syn_tco849 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[13] = 1.825"
syn_tco850 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[14] = 1.806"
syn_tco851 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[15] = 1.752"
syn_tco852 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[16] = 1.743"
syn_tco853 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[17] = 1.775"
syn_tco854 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[18] = 1.753"
syn_tco855 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[19] = 1.722"
syn_tco856 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[20] = 1.787"
syn_tco857 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[21] = 1.811"
syn_tco858 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[22] = 1.737"
syn_tco859 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[23] = 1.796"
syn_tco860 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[24] = 1.768"
syn_tco861 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[25] = 1.768"
syn_tco862 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[26] = 1.762"
syn_tco863 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[27] = 1.796"
syn_tco864 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[28] = 1.793"
syn_tco865 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[2] = 1.739"
syn_tco866 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[3] = 1.728"
syn_tco867 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[4] = 1.744"
syn_tco868 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[5] = 1.731"
syn_tco869 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[6] = 1.855"
syn_tco870 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[7] = 1.822"
syn_tco871 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[8] = 1.763"
syn_tco872 = " FIC_3_PCLK->FIC_3_APB_M_PADDR[9] = 1.716"
syn_tco873 = " FIC_3_PCLK->FIC_3_APB_M_PENABLE = 1.693"
syn_tco874 = " FIC_3_PCLK->FIC_3_APB_M_PSEL = 1.678"
syn_tco875 = " FIC_3_PCLK->FIC_3_APB_M_PSTRB[0] = 1.659"
syn_tco876 = " FIC_3_PCLK->FIC_3_APB_M_PSTRB[1] = 1.609"
syn_tco877 = " FIC_3_PCLK->FIC_3_APB_M_PSTRB[2] = 1.619"
syn_tco878 = " FIC_3_PCLK->FIC_3_APB_M_PSTRB[3] = 1.631"
syn_tco879 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[0] = 1.436"
syn_tco880 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[10] = 1.451"
syn_tco881 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[11] = 1.430"
syn_tco882 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[12] = 1.438"
syn_tco883 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[13] = 1.463"
syn_tco884 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[14] = 1.452"
syn_tco885 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[15] = 1.444"
syn_tco886 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[16] = 1.443"
syn_tco887 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[17] = 1.450"
syn_tco888 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[18] = 1.427"
syn_tco889 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[19] = 1.463"
syn_tco890 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[1] = 1.442"
syn_tco891 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[20] = 1.430"
syn_tco892 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[21] = 1.593"
syn_tco893 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[22] = 1.743"
syn_tco894 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[23] = 1.743"
syn_tco895 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[24] = 1.696"
syn_tco896 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[25] = 1.751"
syn_tco897 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[26] = 1.668"
syn_tco898 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[27] = 1.738"
syn_tco899 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[28] = 1.655"
syn_tco900 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[29] = 1.723"
syn_tco901 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[2] = 1.438"
syn_tco902 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[30] = 1.663"
syn_tco903 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[31] = 1.676"
syn_tco904 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[3] = 1.430"
syn_tco905 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[4] = 1.436"
syn_tco906 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[5] = 1.435"
syn_tco907 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[6] = 1.438"
syn_tco908 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[7] = 1.441"
syn_tco909 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[8] = 1.419"
syn_tco910 = " FIC_3_PCLK->FIC_3_APB_M_PWDATA[9] = 1.443"
syn_tco911 = " FIC_3_PCLK->FIC_3_APB_M_PWRITE = 1.380"
syn_tco912 = " JTAG_TCK_F2M->JTAG_TDO_M2F = 5.484"
syn_tco913 = " JTAG_TCK_F2M->JTAG_TDO_OE_M2F = 5.566"
syn_tco914 = " JTAG_TCK_F2M->JTAG_TDO_M2F = 5.350"
syn_tco915 = " JTAG_TCK_F2M->JTAG_TDO_OE_M2F = 5.474"
syn_tco916 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[0] = 4.653"
syn_tco917 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[100] = 4.352"
syn_tco918 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[101] = 4.021"
syn_tco919 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[102] = 4.149"
syn_tco920 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[103] = 4.129"
syn_tco921 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[104] = 4.316"
syn_tco922 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[105] = 3.914"
syn_tco923 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[106] = 3.939"
syn_tco924 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[107] = 4.137"
syn_tco925 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[108] = 4.023"
syn_tco926 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[109] = 4.164"
syn_tco927 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[10] = 4.564"
syn_tco928 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[110] = 4.208"
syn_tco929 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[111] = 4.233"
syn_tco930 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[112] = 4.241"
syn_tco931 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[113] = 4.446"
syn_tco932 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[114] = 4.192"
syn_tco933 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[115] = 4.140"
syn_tco934 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[116] = 4.213"
syn_tco935 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[117] = 3.820"
syn_tco936 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[118] = 4.262"
syn_tco937 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[119] = 4.202"
syn_tco938 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[11] = 4.742"
syn_tco939 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[120] = 4.401"
syn_tco940 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[121] = 4.194"
syn_tco941 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[122] = 4.315"
syn_tco942 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[123] = 4.434"
syn_tco943 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[124] = 4.555"
syn_tco944 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[125] = 4.333"
syn_tco945 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[126] = 4.310"
syn_tco946 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[127] = 3.998"
syn_tco947 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[12] = 4.645"
syn_tco948 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[13] = 4.662"
syn_tco949 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[14] = 4.639"
syn_tco950 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[15] = 4.613"
syn_tco951 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[16] = 4.475"
syn_tco952 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[17] = 4.458"
syn_tco953 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[18] = 4.386"
syn_tco954 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[19] = 4.505"
syn_tco955 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[1] = 4.688"
syn_tco956 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[20] = 4.396"
syn_tco957 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[21] = 4.568"
syn_tco958 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[22] = 4.462"
syn_tco959 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[23] = 4.474"
syn_tco960 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[24] = 4.394"
syn_tco961 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[25] = 4.380"
syn_tco962 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[26] = 4.482"
syn_tco963 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[27] = 4.306"
syn_tco964 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[28] = 4.275"
syn_tco965 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[29] = 4.327"
syn_tco966 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[2] = 4.694"
syn_tco967 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[30] = 4.462"
syn_tco968 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[31] = 4.344"
syn_tco969 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[32] = 4.376"
syn_tco970 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[33] = 4.468"
syn_tco971 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[34] = 4.474"
syn_tco972 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[35] = 4.382"
syn_tco973 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[36] = 4.293"
syn_tco974 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[37] = 4.335"
syn_tco975 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[38] = 4.218"
syn_tco976 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[39] = 4.290"
syn_tco977 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[3] = 4.723"
syn_tco978 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[40] = 4.267"
syn_tco979 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[41] = 4.372"
syn_tco980 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[42] = 4.431"
syn_tco981 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[43] = 4.448"
syn_tco982 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[44] = 4.411"
syn_tco983 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[45] = 4.438"
syn_tco984 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[46] = 4.538"
syn_tco985 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[47] = 4.353"
syn_tco986 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[48] = 4.245"
syn_tco987 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[49] = 4.326"
syn_tco988 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[4] = 4.610"
syn_tco989 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[50] = 4.266"
syn_tco990 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[51] = 4.099"
syn_tco991 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[52] = 4.161"
syn_tco992 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[53] = 4.075"
syn_tco993 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[54] = 4.111"
syn_tco994 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[55] = 4.036"
syn_tco995 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[56] = 4.085"
syn_tco996 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[57] = 4.002"
syn_tco997 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[58] = 4.018"
syn_tco998 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[59] = 4.173"
syn_tco999 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[5] = 4.650"
syn_tco1000 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[60] = 4.144"
syn_tco1001 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[61] = 4.206"
syn_tco1002 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[62] = 4.153"
syn_tco1003 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[63] = 4.377"
syn_tco1004 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[64] = 4.242"
syn_tco1005 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[65] = 4.211"
syn_tco1006 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[66] = 4.237"
syn_tco1007 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[67] = 4.211"
syn_tco1008 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[68] = 4.343"
syn_tco1009 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[69] = 4.045"
syn_tco1010 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[6] = 4.570"
syn_tco1011 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[70] = 4.392"
syn_tco1012 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[71] = 4.378"
syn_tco1013 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[72] = 4.163"
syn_tco1014 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[73] = 4.212"
syn_tco1015 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[74] = 4.263"
syn_tco1016 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[75] = 4.295"
syn_tco1017 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[76] = 4.220"
syn_tco1018 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[77] = 4.462"
syn_tco1019 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[78] = 4.306"
syn_tco1020 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[79] = 4.290"
syn_tco1021 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[7] = 4.680"
syn_tco1022 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[80] = 4.375"
syn_tco1023 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[81] = 4.342"
syn_tco1024 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[82] = 4.371"
syn_tco1025 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[83] = 4.231"
syn_tco1026 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[84] = 4.208"
syn_tco1027 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[85] = 4.347"
syn_tco1028 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[86] = 4.030"
syn_tco1029 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[87] = 4.120"
syn_tco1030 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[88] = 4.101"
syn_tco1031 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[89] = 4.297"
syn_tco1032 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[8] = 4.682"
syn_tco1033 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[90] = 4.124"
syn_tco1034 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[91] = 4.335"
syn_tco1035 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[92] = 4.360"
syn_tco1036 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[93] = 4.223"
syn_tco1037 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[94] = 4.195"
syn_tco1038 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[95] = 4.150"
syn_tco1039 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[96] = 4.181"
syn_tco1040 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[97] = 4.042"
syn_tco1041 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[98] = 4.172"
syn_tco1042 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[99] = 4.015"
syn_tco1043 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DATA_M2F[9] = 4.667"
syn_tco1044 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DA_STB_M2F = 2.985"
syn_tco1045 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_DP_STB_M2F = 3.303"
syn_tco1046 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_IPV6_M2F = 3.136"
syn_tco1047 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_IP_DA_STB_M2F = 3.260"
syn_tco1048 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_IP_SA_STB_M2F = 3.241"
syn_tco1049 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_SA_STB_M2F = 3.161"
syn_tco1050 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_SP_STB_M2F = 3.141"
syn_tco1051 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_TYPE_STB_M2F = 3.169"
syn_tco1052 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_VLAN_TAG1_STB_M2F = 3.123"
syn_tco1053 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_FILTER_VLAN_TAG2_STB_M2F = 3.223"
syn_tco1054 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_TSU_DELAY_REQ_RX_M2F = 3.673"
syn_tco1055 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_TSU_PDELAY_REQ_RX_M2F = 3.528"
syn_tco1056 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_TSU_PDELAY_RESP_RX_M2F = 3.498"
syn_tco1057 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_TSU_SOF_RX_M2F = 3.402"
syn_tco1058 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_TSU_SYNC_FRAME_RX_M2F = 3.581"
syn_tco1059 = " MAC_0_GMII_MII_RX_CLK_F2M->MAC_0_WOL_M2F = 3.131"
syn_tco1060 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_GMII_MII_TXD_M2F[0] = 2.501"
syn_tco1061 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_GMII_MII_TXD_M2F[1] = 2.439"
syn_tco1062 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_GMII_MII_TXD_M2F[2] = 2.496"
syn_tco1063 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_GMII_MII_TXD_M2F[3] = 2.445"
syn_tco1064 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_GMII_MII_TXD_M2F[4] = 2.494"
syn_tco1065 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_GMII_MII_TXD_M2F[5] = 2.488"
syn_tco1066 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_GMII_MII_TXD_M2F[6] = 2.460"
syn_tco1067 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_GMII_MII_TXD_M2F[7] = 2.512"
syn_tco1068 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_GMII_MII_TX_EN_M2F = 2.520"
syn_tco1069 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_GMII_MII_TX_ER_M2F = 2.493"
syn_tco1070 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_TSU_DELAY_REQ_TX_M2F = 3.586"
syn_tco1071 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_TSU_PDELAY_REQ_TX_M2F = 3.402"
syn_tco1072 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_TSU_PDELAY_RESP_TX_M2F = 3.235"
syn_tco1073 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_TSU_SOF_TX_M2F = 3.344"
syn_tco1074 = " MAC_0_GMII_MII_TX_CLK_F2M->MAC_0_TSU_SYNC_FRAME_TX_M2F = 3.263"
syn_tco1075 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CMP_VAL_M2F = 2.848"
syn_tco1076 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[0] = 2.985"
syn_tco1077 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[10] = 2.949"
syn_tco1078 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[11] = 2.722"
syn_tco1079 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[12] = 2.912"
syn_tco1080 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[13] = 2.899"
syn_tco1081 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[14] = 2.925"
syn_tco1082 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[15] = 2.879"
syn_tco1083 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[16] = 2.937"
syn_tco1084 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[17] = 2.744"
syn_tco1085 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[18] = 2.769"
syn_tco1086 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[19] = 2.852"
syn_tco1087 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[1] = 2.683"
syn_tco1088 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[20] = 3.117"
syn_tco1089 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[21] = 2.936"
syn_tco1090 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[22] = 2.982"
syn_tco1091 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[23] = 2.844"
syn_tco1092 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[24] = 3.142"
syn_tco1093 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[25] = 2.845"
syn_tco1094 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[26] = 2.788"
syn_tco1095 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[27] = 3.062"
syn_tco1096 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[28] = 2.845"
syn_tco1097 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[29] = 2.737"
syn_tco1098 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[2] = 2.709"
syn_tco1099 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[30] = 3.028"
syn_tco1100 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[31] = 2.878"
syn_tco1101 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[32] = 2.924"
syn_tco1102 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[33] = 3.003"
syn_tco1103 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[34] = 2.869"
syn_tco1104 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[35] = 2.994"
syn_tco1105 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[36] = 2.958"
syn_tco1106 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[37] = 2.953"
syn_tco1107 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[38] = 2.836"
syn_tco1108 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[39] = 3.172"
syn_tco1109 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[3] = 2.828"
syn_tco1110 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[40] = 2.769"
syn_tco1111 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[41] = 3.044"
syn_tco1112 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[42] = 2.807"
syn_tco1113 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[43] = 3.060"
syn_tco1114 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[44] = 3.032"
syn_tco1115 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[45] = 2.901"
syn_tco1116 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[46] = 2.986"
syn_tco1117 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[47] = 3.130"
syn_tco1118 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[48] = 2.907"
syn_tco1119 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[49] = 2.834"
syn_tco1120 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[4] = 2.677"
syn_tco1121 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[50] = 3.143"
syn_tco1122 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[51] = 3.091"
syn_tco1123 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[52] = 2.978"
syn_tco1124 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[53] = 2.918"
syn_tco1125 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[54] = 3.098"
syn_tco1126 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[55] = 2.994"
syn_tco1127 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[56] = 3.104"
syn_tco1128 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[57] = 2.982"
syn_tco1129 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[58] = 3.069"
syn_tco1130 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[59] = 2.893"
syn_tco1131 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[5] = 3.030"
syn_tco1132 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[60] = 3.108"
syn_tco1133 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[61] = 2.907"
syn_tco1134 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[62] = 2.827"
syn_tco1135 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[63] = 2.823"
syn_tco1136 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[64] = 2.917"
syn_tco1137 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[65] = 2.894"
syn_tco1138 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[66] = 2.894"
syn_tco1139 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[67] = 2.958"
syn_tco1140 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[68] = 2.920"
syn_tco1141 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[69] = 2.906"
syn_tco1142 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[6] = 2.919"
syn_tco1143 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[70] = 2.900"
syn_tco1144 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[71] = 2.869"
syn_tco1145 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[72] = 3.141"
syn_tco1146 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[73] = 2.780"
syn_tco1147 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[74] = 2.825"
syn_tco1148 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[75] = 2.813"
syn_tco1149 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[76] = 2.948"
syn_tco1150 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[77] = 2.878"
syn_tco1151 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[78] = 2.763"
syn_tco1152 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[79] = 2.878"
syn_tco1153 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[7] = 2.922"
syn_tco1154 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[80] = 2.785"
syn_tco1155 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[81] = 2.771"
syn_tco1156 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[82] = 2.989"
syn_tco1157 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[83] = 2.711"
syn_tco1158 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[84] = 2.801"
syn_tco1159 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[85] = 2.974"
syn_tco1160 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[86] = 2.943"
syn_tco1161 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[87] = 3.021"
syn_tco1162 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[88] = 2.870"
syn_tco1163 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[89] = 2.869"
syn_tco1164 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[8] = 2.869"
syn_tco1165 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[90] = 3.049"
syn_tco1166 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[91] = 2.921"
syn_tco1167 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[92] = 2.964"
syn_tco1168 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[93] = 2.944"
syn_tco1169 = " MAC_0_TSU_CLK_F2M->MAC_0_TSU_TIMER_CNT_M2F[9] = 2.869"
syn_tco1170 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[0] = 5.038"
syn_tco1171 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[100] = 4.631"
syn_tco1172 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[101] = 4.723"
syn_tco1173 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[102] = 4.643"
syn_tco1174 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[103] = 4.642"
syn_tco1175 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[104] = 4.772"
syn_tco1176 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[105] = 4.685"
syn_tco1177 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[106] = 4.772"
syn_tco1178 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[107] = 4.719"
syn_tco1179 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[108] = 4.675"
syn_tco1180 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[109] = 4.685"
syn_tco1181 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[10] = 4.889"
syn_tco1182 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[110] = 4.745"
syn_tco1183 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[111] = 4.698"
syn_tco1184 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[112] = 4.590"
syn_tco1185 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[113] = 4.737"
syn_tco1186 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[114] = 4.578"
syn_tco1187 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[115] = 4.729"
syn_tco1188 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[116] = 4.651"
syn_tco1189 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[117] = 4.726"
syn_tco1190 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[118] = 4.734"
syn_tco1191 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[119] = 4.532"
syn_tco1192 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[11] = 4.999"
syn_tco1193 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[120] = 4.635"
syn_tco1194 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[121] = 4.662"
syn_tco1195 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[122] = 4.694"
syn_tco1196 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[123] = 4.623"
syn_tco1197 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[124] = 4.710"
syn_tco1198 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[125] = 4.607"
syn_tco1199 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[126] = 4.699"
syn_tco1200 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[127] = 4.660"
syn_tco1201 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[12] = 5.050"
syn_tco1202 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[13] = 4.838"
syn_tco1203 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[14] = 4.836"
syn_tco1204 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[15] = 4.967"
syn_tco1205 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[16] = 4.895"
syn_tco1206 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[17] = 4.856"
syn_tco1207 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[18] = 5.044"
syn_tco1208 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[19] = 4.904"
syn_tco1209 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[1] = 4.882"
syn_tco1210 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[20] = 4.910"
syn_tco1211 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[21] = 4.847"
syn_tco1212 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[22] = 4.788"
syn_tco1213 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[23] = 4.968"
syn_tco1214 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[24] = 4.782"
syn_tco1215 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[25] = 5.010"
syn_tco1216 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[26] = 4.845"
syn_tco1217 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[27] = 4.844"
syn_tco1218 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[28] = 4.929"
syn_tco1219 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[29] = 4.884"
syn_tco1220 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[2] = 4.933"
syn_tco1221 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[30] = 4.826"
syn_tco1222 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[31] = 4.645"
syn_tco1223 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[32] = 4.722"
syn_tco1224 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[33] = 4.772"
syn_tco1225 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[34] = 4.537"
syn_tco1226 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[35] = 4.769"
syn_tco1227 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[36] = 4.695"
syn_tco1228 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[37] = 4.609"
syn_tco1229 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[38] = 4.757"
syn_tco1230 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[39] = 4.760"
syn_tco1231 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[3] = 5.179"
syn_tco1232 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[40] = 4.637"
syn_tco1233 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[41] = 4.620"
syn_tco1234 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[42] = 4.684"
syn_tco1235 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[43] = 4.600"
syn_tco1236 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[44] = 4.640"
syn_tco1237 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[45] = 4.637"
syn_tco1238 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[46] = 4.676"
syn_tco1239 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[47] = 4.710"
syn_tco1240 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[48] = 4.758"
syn_tco1241 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[49] = 4.652"
syn_tco1242 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[4] = 4.986"
syn_tco1243 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[50] = 4.745"
syn_tco1244 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[51] = 4.635"
syn_tco1245 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[52] = 4.747"
syn_tco1246 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[53] = 4.627"
syn_tco1247 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[54] = 4.739"
syn_tco1248 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[55] = 4.693"
syn_tco1249 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[56] = 4.680"
syn_tco1250 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[57] = 4.678"
syn_tco1251 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[58] = 4.615"
syn_tco1252 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[59] = 4.608"
syn_tco1253 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[5] = 4.831"
syn_tco1254 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[60] = 4.695"
syn_tco1255 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[61] = 4.694"
syn_tco1256 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[62] = 4.651"
syn_tco1257 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[63] = 4.691"
syn_tco1258 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[64] = 4.816"
syn_tco1259 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[65] = 4.741"
syn_tco1260 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[66] = 4.730"
syn_tco1261 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[67] = 4.814"
syn_tco1262 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[68] = 4.599"
syn_tco1263 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[69] = 4.722"
syn_tco1264 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[6] = 4.971"
syn_tco1265 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[70] = 4.722"
syn_tco1266 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[71] = 4.799"
syn_tco1267 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[72] = 4.828"
syn_tco1268 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[73] = 4.713"
syn_tco1269 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[74] = 4.550"
syn_tco1270 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[75] = 4.639"
syn_tco1271 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[76] = 4.672"
syn_tco1272 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[77] = 4.622"
syn_tco1273 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[78] = 4.615"
syn_tco1274 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[79] = 4.702"
syn_tco1275 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[7] = 4.811"
syn_tco1276 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[80] = 4.654"
syn_tco1277 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[81] = 4.677"
syn_tco1278 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[82] = 4.624"
syn_tco1279 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[83] = 4.691"
syn_tco1280 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[84] = 4.811"
syn_tco1281 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[85] = 4.623"
syn_tco1282 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[86] = 4.684"
syn_tco1283 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[87] = 4.622"
syn_tco1284 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[88] = 4.624"
syn_tco1285 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[89] = 4.719"
syn_tco1286 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[8] = 4.873"
syn_tco1287 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[90] = 4.662"
syn_tco1288 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[91] = 4.706"
syn_tco1289 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[92] = 4.683"
syn_tco1290 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[93] = 4.690"
syn_tco1291 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[94] = 4.584"
syn_tco1292 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[95] = 4.585"
syn_tco1293 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[96] = 4.774"
syn_tco1294 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[97] = 4.870"
syn_tco1295 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[98] = 4.771"
syn_tco1296 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[99] = 4.724"
syn_tco1297 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DATA_M2F[9] = 4.977"
syn_tco1298 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DA_STB_M2F = 3.607"
syn_tco1299 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_DP_STB_M2F = 3.695"
syn_tco1300 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_IPV6_M2F = 3.521"
syn_tco1301 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_IP_DA_STB_M2F = 3.553"
syn_tco1302 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_IP_SA_STB_M2F = 3.481"
syn_tco1303 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_SA_STB_M2F = 3.491"
syn_tco1304 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_SP_STB_M2F = 3.536"
syn_tco1305 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_TYPE_STB_M2F = 3.508"
syn_tco1306 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_VLAN_TAG1_STB_M2F = 3.550"
syn_tco1307 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_FILTER_VLAN_TAG2_STB_M2F = 3.564"
syn_tco1308 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_TSU_DELAY_REQ_RX_M2F = 3.993"
syn_tco1309 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_TSU_PDELAY_REQ_RX_M2F = 3.697"
syn_tco1310 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_TSU_PDELAY_RESP_RX_M2F = 3.744"
syn_tco1311 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_TSU_SOF_RX_M2F = 3.799"
syn_tco1312 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_TSU_SYNC_FRAME_RX_M2F = 4.021"
syn_tco1313 = " MAC_1_GMII_MII_RX_CLK_F2M->MAC_1_WOL_M2F = 3.435"
syn_tco1314 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_GMII_MII_TXD_M2F[0] = 2.711"
syn_tco1315 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_GMII_MII_TXD_M2F[1] = 2.636"
syn_tco1316 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_GMII_MII_TXD_M2F[2] = 2.639"
syn_tco1317 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_GMII_MII_TXD_M2F[3] = 2.662"
syn_tco1318 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_GMII_MII_TXD_M2F[4] = 2.672"
syn_tco1319 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_GMII_MII_TXD_M2F[5] = 2.631"
syn_tco1320 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_GMII_MII_TXD_M2F[6] = 2.642"
syn_tco1321 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_GMII_MII_TXD_M2F[7] = 2.645"
syn_tco1322 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_GMII_MII_TX_EN_M2F = 2.615"
syn_tco1323 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_GMII_MII_TX_ER_M2F = 2.612"
syn_tco1324 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_TSU_DELAY_REQ_TX_M2F = 3.901"
syn_tco1325 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_TSU_PDELAY_REQ_TX_M2F = 3.753"
syn_tco1326 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_TSU_PDELAY_RESP_TX_M2F = 3.789"
syn_tco1327 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_TSU_SOF_TX_M2F = 3.641"
syn_tco1328 = " MAC_1_GMII_MII_TX_CLK_F2M->MAC_1_TSU_SYNC_FRAME_TX_M2F = 3.651"
syn_tco1329 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CMP_VAL_M2F = 3.902"
syn_tco1330 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[0] = 3.725"
syn_tco1331 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[10] = 3.689"
syn_tco1332 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[11] = 3.734"
syn_tco1333 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[12] = 3.638"
syn_tco1334 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[13] = 3.793"
syn_tco1335 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[14] = 3.668"
syn_tco1336 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[15] = 3.728"
syn_tco1337 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[16] = 3.680"
syn_tco1338 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[17] = 3.607"
syn_tco1339 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[18] = 3.775"
syn_tco1340 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[19] = 3.528"
syn_tco1341 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[1] = 3.799"
syn_tco1342 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[20] = 3.722"
syn_tco1343 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[21] = 3.865"
syn_tco1344 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[22] = 3.684"
syn_tco1345 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[23] = 3.740"
syn_tco1346 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[24] = 3.620"
syn_tco1347 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[25] = 3.745"
syn_tco1348 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[26] = 3.678"
syn_tco1349 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[27] = 3.606"
syn_tco1350 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[28] = 3.538"
syn_tco1351 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[29] = 3.674"
syn_tco1352 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[2] = 3.752"
syn_tco1353 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[30] = 3.823"
syn_tco1354 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[31] = 3.681"
syn_tco1355 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[32] = 3.808"
syn_tco1356 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[33] = 3.725"
syn_tco1357 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[34] = 3.808"
syn_tco1358 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[35] = 3.828"
syn_tco1359 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[36] = 3.868"
syn_tco1360 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[37] = 3.759"
syn_tco1361 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[38] = 3.878"
syn_tco1362 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[39] = 3.768"
syn_tco1363 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[3] = 3.739"
syn_tco1364 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[40] = 3.915"
syn_tco1365 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[41] = 3.653"
syn_tco1366 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[42] = 3.542"
syn_tco1367 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[43] = 3.766"
syn_tco1368 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[44] = 3.727"
syn_tco1369 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[45] = 3.908"
syn_tco1370 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[46] = 3.714"
syn_tco1371 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[47] = 3.555"
syn_tco1372 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[48] = 3.465"
syn_tco1373 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[49] = 3.619"
syn_tco1374 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[4] = 3.704"
syn_tco1375 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[50] = 3.829"
syn_tco1376 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[51] = 3.632"
syn_tco1377 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[52] = 3.599"
syn_tco1378 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[53] = 3.664"
syn_tco1379 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[54] = 3.637"
syn_tco1380 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[55] = 3.621"
syn_tco1381 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[56] = 3.687"
syn_tco1382 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[57] = 3.731"
syn_tco1383 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[58] = 3.560"
syn_tco1384 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[59] = 3.578"
syn_tco1385 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[5] = 3.758"
syn_tco1386 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[60] = 3.490"
syn_tco1387 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[61] = 3.591"
syn_tco1388 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[62] = 3.583"
syn_tco1389 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[63] = 3.712"
syn_tco1390 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[64] = 3.635"
syn_tco1391 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[65] = 3.497"
syn_tco1392 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[66] = 3.644"
syn_tco1393 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[67] = 3.727"
syn_tco1394 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[68] = 3.599"
syn_tco1395 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[69] = 3.776"
syn_tco1396 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[6] = 3.766"
syn_tco1397 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[70] = 3.672"
syn_tco1398 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[71] = 3.717"
syn_tco1399 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[72] = 3.655"
syn_tco1400 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[73] = 3.709"
syn_tco1401 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[74] = 3.735"
syn_tco1402 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[75] = 3.661"
syn_tco1403 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[76] = 3.468"
syn_tco1404 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[77] = 3.752"
syn_tco1405 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[78] = 3.744"
syn_tco1406 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[79] = 3.644"
syn_tco1407 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[7] = 3.735"
syn_tco1408 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[80] = 3.481"
syn_tco1409 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[81] = 3.575"
syn_tco1410 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[82] = 3.622"
syn_tco1411 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[83] = 3.463"
syn_tco1412 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[84] = 3.767"
syn_tco1413 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[85] = 3.561"
syn_tco1414 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[86] = 3.637"
syn_tco1415 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[87] = 3.740"
syn_tco1416 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[88] = 3.838"
syn_tco1417 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[89] = 3.885"
syn_tco1418 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[8] = 3.818"
syn_tco1419 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[90] = 3.882"
syn_tco1420 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[91] = 3.802"
syn_tco1421 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[92] = 3.814"
syn_tco1422 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[93] = 3.911"
syn_tco1423 = " MAC_1_TSU_CLK_F2M->MAC_1_TSU_TIMER_CNT_M2F[9] = 3.904"
syn_tpd1424 = " SPARE_1_F2M[0]->MSSIO0_OUT = 4.368"
syn_tpd1425 = " SPARE_1_F2M[10]->MSSIO10_OUT = 3.754"
syn_tpd1426 = " SPARE_1_F2M[11]->MSSIO11_OUT = 3.620"
syn_tpd1427 = " SPARE_1_F2M[12]->MSSIO12_OUT = 3.550"
syn_tpd1428 = " SPARE_1_F2M[13]->MSSIO13_OUT = 3.854"
syn_tpd1429 = " SPARE_1_F2M[14]->MSSIO14_OUT = 4.039"
syn_tpd1430 = " SPARE_1_F2M[15]->MSSIO15_OUT = 3.605"
syn_tpd1431 = " SPARE_1_F2M[16]->MSSIO16_OUT = 3.519"
syn_tpd1432 = " SPARE_1_F2M[17]->MSSIO17_OUT = 3.630"
syn_tpd1433 = " SPARE_1_F2M[18]->MSSIO18_OUT = 3.359"
syn_tpd1434 = " SPARE_1_F2M[19]->MSSIO19_OUT = 3.351"
syn_tpd1435 = " SPARE_1_F2M[1]->MSSIO1_OUT = 4.249"
syn_tpd1436 = " SPARE_1_F2M[20]->MSSIO20_OUT = 3.625"
syn_tpd1437 = " SPARE_1_F2M[21]->MSSIO21_OUT = 3.419"
syn_tpd1438 = " SPARE_1_F2M[22]->MSSIO22_OUT = 3.489"
syn_tpd1439 = " SPARE_1_F2M[23]->MSSIO23_OUT = 3.848"
syn_tpd1440 = " SPARE_1_F2M[24]->MSSIO24_OUT = 3.671"
syn_tpd1441 = " SPARE_1_F2M[25]->MSSIO25_OUT = 3.845"
syn_tpd1442 = " SPARE_1_F2M[26]->MSSIO26_OUT = 3.683"
syn_tpd1443 = " SPARE_1_F2M[27]->MSSIO27_OUT = 3.619"
syn_tpd1444 = " SPARE_1_F2M[28]->MSSIO28_OUT = 3.538"
syn_tpd1445 = " SPARE_1_F2M[29]->MSSIO29_OUT = 3.637"
syn_tpd1446 = " SPARE_1_F2M[2]->MSSIO2_OUT = 3.998"
syn_tpd1447 = " SPARE_1_F2M[30]->MSSIO30_OUT = 4.223"
syn_tpd1448 = " SPARE_1_F2M[31]->MSSIO31_OUT = 3.978"
syn_tpd1449 = " SPARE_1_F2M[32]->MSSIO32_OUT = 3.596"
syn_tpd1450 = " SPARE_1_F2M[33]->MSSIO33_OUT = 3.679"
syn_tpd1451 = " SPARE_1_F2M[34]->MSSIO34_OUT = 3.334"
syn_tpd1452 = " SPARE_1_F2M[35]->MSSIO35_OUT = 3.758"
syn_tpd1453 = " SPARE_1_F2M[36]->MSSIO36_OUT = 3.747"
syn_tpd1454 = " SPARE_1_F2M[37]->MSSIO37_OUT = 3.903"
syn_tpd1455 = " SPARE_1_F2M[3]->MSSIO3_OUT = 3.822"
syn_tpd1456 = " SPARE_1_F2M[4]->MSSIO4_OUT = 4.228"
syn_tpd1457 = " SPARE_1_F2M[5]->MSSIO5_OUT = 4.322"
syn_tpd1458 = " SPARE_1_F2M[6]->MSSIO6_OUT = 4.203"
syn_tpd1459 = " SPARE_1_F2M[7]->MSSIO7_OUT = 3.627"
syn_tpd1460 = " SPARE_1_F2M[8]->MSSIO8_OUT = 3.611"
syn_tpd1461 = " SPARE_1_F2M[9]->MSSIO9_OUT = 3.813"
syn_tpd1462 = " SPARE_2_F2M[0]->MSSIO0_OE = 4.555"
syn_tpd1463 = " SPARE_2_F2M[10]->MSSIO10_OE = 3.567"
syn_tpd1464 = " SPARE_2_F2M[11]->MSSIO11_OE = 4.497"
syn_tpd1465 = " SPARE_2_F2M[12]->MSSIO12_OE = 3.346"
syn_tpd1466 = " SPARE_2_F2M[13]->MSSIO13_OE = 4.265"
syn_tpd1467 = " SPARE_2_F2M[14]->MSSIO14_OE = 3.749"
syn_tpd1468 = " SPARE_2_F2M[15]->MSSIO15_OE = 4.143"
syn_tpd1469 = " SPARE_2_F2M[16]->MSSIO16_OE = 3.511"
syn_tpd1470 = " SPARE_2_F2M[17]->MSSIO17_OE = 3.843"
syn_tpd1471 = " SPARE_2_F2M[18]->MSSIO18_OE = 3.423"
syn_tpd1472 = " SPARE_2_F2M[19]->MSSIO19_OE = 3.643"
syn_tpd1473 = " SPARE_2_F2M[1]->MSSIO1_OE = 4.140"
syn_tpd1474 = " SPARE_2_F2M[20]->MSSIO20_OE = 3.400"
syn_tpd1475 = " SPARE_2_F2M[21]->MSSIO21_OE = 3.380"
syn_tpd1476 = " SPARE_2_F2M[22]->MSSIO22_OE = 3.766"
syn_tpd1477 = " SPARE_2_F2M[23]->MSSIO23_OE = 4.617"
syn_tpd1478 = " SPARE_2_F2M[24]->MSSIO24_OE = 3.832"
syn_tpd1479 = " SPARE_2_F2M[25]->MSSIO25_OE = 3.730"
syn_tpd1480 = " SPARE_2_F2M[26]->MSSIO26_OE = 4.001"
syn_tpd1481 = " SPARE_2_F2M[27]->MSSIO27_OE = 3.873"
syn_tpd1482 = " SPARE_2_F2M[28]->MSSIO28_OE = 4.261"
syn_tpd1483 = " SPARE_2_F2M[29]->MSSIO29_OE = 3.583"
syn_tpd1484 = " SPARE_2_F2M[2]->MSSIO2_OE = 3.995"
syn_tpd1485 = " SPARE_2_F2M[30]->MSSIO30_OE = 4.527"
syn_tpd1486 = " SPARE_2_F2M[31]->MSSIO31_OE = 4.356"
syn_tpd1487 = " SPARE_2_F2M[32]->MSSIO32_OE = 4.177"
syn_tpd1488 = " SPARE_2_F2M[33]->MSSIO33_OE = 4.136"
syn_tpd1489 = " SPARE_2_F2M[34]->MSSIO34_OE = 4.069"
syn_tpd1490 = " SPARE_2_F2M[35]->MSSIO35_OE = 3.701"
syn_tpd1491 = " SPARE_2_F2M[36]->MSSIO36_OE = 4.030"
syn_tpd1492 = " SPARE_2_F2M[37]->MSSIO37_OE = 4.514"
syn_tpd1493 = " SPARE_2_F2M[3]->MSSIO3_OE = 4.127"
syn_tpd1494 = " SPARE_2_F2M[4]->MSSIO4_OE = 4.173"
syn_tpd1495 = " SPARE_2_F2M[5]->MSSIO5_OE = 4.348"
syn_tpd1496 = " SPARE_2_F2M[6]->MSSIO6_OE = 4.196"
syn_tpd1497 = " SPARE_2_F2M[7]->MSSIO7_OE = 3.790"
syn_tpd1498 = " SPARE_2_F2M[8]->MSSIO8_OE = 3.582"
syn_tpd1499 = " SPARE_2_F2M[9]->MSSIO9_OE = 4.427"
syn_tpd1500 = " SPI_0_SS_F2M->SPI_0_DO_OE_M2F = 2.254"
syn_tpd1501 = " SPI_1_SS_F2M->SPI_1_DO_OE_M2F = 3.008"
*/
/* synthesis black_box_pad_pin ="" */
input  FIC_0_ACLK;
input  FIC_0_AXI4_M_AWREADY;
input  FIC_0_AXI4_M_WREADY;
input  [7:0] FIC_0_AXI4_M_BID;
input  [1:0] FIC_0_AXI4_M_BRESP;
input  FIC_0_AXI4_M_BVALID;
input  FIC_0_AXI4_M_ARREADY;
input  [7:0] FIC_0_AXI4_M_RID;
input  [63:0] FIC_0_AXI4_M_RDATA;
input  [1:0] FIC_0_AXI4_M_RRESP;
input  FIC_0_AXI4_M_RLAST;
input  FIC_0_AXI4_M_RVALID;
input  [3:0] FIC_0_AXI4_S_AWID;
input  [37:0] FIC_0_AXI4_S_AWADDR;
input  [7:0] FIC_0_AXI4_S_AWLEN;
input  [2:0] FIC_0_AXI4_S_AWSIZE;
input  [1:0] FIC_0_AXI4_S_AWBURST;
input  [3:0] FIC_0_AXI4_S_AWQOS;
input  FIC_0_AXI4_S_AWLOCK;
input  [3:0] FIC_0_AXI4_S_AWCACHE;
input  [2:0] FIC_0_AXI4_S_AWPROT;
input  FIC_0_AXI4_S_AWVALID;
input  [63:0] FIC_0_AXI4_S_WDATA;
input  [7:0] FIC_0_AXI4_S_WSTRB;
input  FIC_0_AXI4_S_WLAST;
input  FIC_0_AXI4_S_WVALID;
input  FIC_0_AXI4_S_BREADY;
input  [3:0] FIC_0_AXI4_S_ARID;
input  [37:0] FIC_0_AXI4_S_ARADDR;
input  [7:0] FIC_0_AXI4_S_ARLEN;
input  [2:0] FIC_0_AXI4_S_ARSIZE;
input  [1:0] FIC_0_AXI4_S_ARBURST;
input  [3:0] FIC_0_AXI4_S_ARQOS;
input  FIC_0_AXI4_S_ARLOCK;
input  [3:0] FIC_0_AXI4_S_ARCACHE;
input  [2:0] FIC_0_AXI4_S_ARPROT;
input  FIC_0_AXI4_S_ARVALID;
input  FIC_0_AXI4_S_RREADY;
input  FIC_1_ACLK;
input  FIC_1_AXI4_M_AWREADY;
input  FIC_1_AXI4_M_WREADY;
input  [7:0] FIC_1_AXI4_M_BID;
input  [1:0] FIC_1_AXI4_M_BRESP;
input  FIC_1_AXI4_M_BVALID;
input  FIC_1_AXI4_M_ARREADY;
input  [7:0] FIC_1_AXI4_M_RID;
input  [63:0] FIC_1_AXI4_M_RDATA;
input  [1:0] FIC_1_AXI4_M_RRESP;
input  FIC_1_AXI4_M_RLAST;
input  FIC_1_AXI4_M_RVALID;
input  [3:0] FIC_1_AXI4_S_AWID;
input  [37:0] FIC_1_AXI4_S_AWADDR;
input  [7:0] FIC_1_AXI4_S_AWLEN;
input  [2:0] FIC_1_AXI4_S_AWSIZE;
input  [1:0] FIC_1_AXI4_S_AWBURST;
input  FIC_1_AXI4_S_AWLOCK;
input  [3:0] FIC_1_AXI4_S_AWCACHE;
input  [3:0] FIC_1_AXI4_S_AWQOS;
input  [2:0] FIC_1_AXI4_S_AWPROT;
input  FIC_1_AXI4_S_AWVALID;
input  [63:0] FIC_1_AXI4_S_WDATA;
input  [7:0] FIC_1_AXI4_S_WSTRB;
input  FIC_1_AXI4_S_WLAST;
input  FIC_1_AXI4_S_WVALID;
input  FIC_1_AXI4_S_BREADY;
input  [3:0] FIC_1_AXI4_S_ARID;
input  [37:0] FIC_1_AXI4_S_ARADDR;
input  [7:0] FIC_1_AXI4_S_ARLEN;
input  [2:0] FIC_1_AXI4_S_ARSIZE;
input  [1:0] FIC_1_AXI4_S_ARBURST;
input  [3:0] FIC_1_AXI4_S_ARQOS;
input  FIC_1_AXI4_S_ARLOCK;
input  [3:0] FIC_1_AXI4_S_ARCACHE;
input  [2:0] FIC_1_AXI4_S_ARPROT;
input  FIC_1_AXI4_S_ARVALID;
input  FIC_1_AXI4_S_RREADY;
input  FIC_2_ACLK;
input  SPARE_3_F2M;
input  [3:0] FIC_2_AXI4_S_AWID;
input  [37:0] FIC_2_AXI4_S_AWADDR;
input  [7:0] FIC_2_AXI4_S_AWLEN;
input  [2:0] FIC_2_AXI4_S_AWSIZE;
input  [1:0] FIC_2_AXI4_S_AWBURST;
input  FIC_2_AXI4_S_AWLOCK;
input  [3:0] FIC_2_AXI4_S_AWCACHE;
input  [3:0] FIC_2_AXI4_S_AWQOS;
input  [2:0] FIC_2_AXI4_S_AWPROT;
input  FIC_2_AXI4_S_AWVALID;
input  [63:0] FIC_2_AXI4_S_WDATA;
input  [7:0] FIC_2_AXI4_S_WSTRB;
input  FIC_2_AXI4_S_WLAST;
input  FIC_2_AXI4_S_WVALID;
input  FIC_2_AXI4_S_BREADY;
input  [3:0] FIC_2_AXI4_S_ARID;
input  [37:0] FIC_2_AXI4_S_ARADDR;
input  [7:0] FIC_2_AXI4_S_ARLEN;
input  [2:0] FIC_2_AXI4_S_ARSIZE;
input  [1:0] FIC_2_AXI4_S_ARBURST;
input  FIC_2_AXI4_S_ARLOCK;
input  [3:0] FIC_2_AXI4_S_ARCACHE;
input  [3:0] FIC_2_AXI4_S_ARQOS;
input  [2:0] FIC_2_AXI4_S_ARPROT;
input  FIC_2_AXI4_S_ARVALID;
input  FIC_2_AXI4_S_RREADY;
input  FIC_3_PCLK;
input  SPARE_4_F2M;
input  [31:0] FIC_3_APB_M_PRDATA;
input  FIC_3_APB_M_PREADY;
input  FIC_3_APB_M_PSLVERR;
input  MMUART_0_DCD_F2M;
input  MMUART_0_RI_F2M;
input  MMUART_0_DSR_F2M;
input  MMUART_0_CTS_F2M;
input  MMUART_0_RXD_F2M;
input  MMUART_0_CLK_F2M;
input  MMUART_1_DCD_F2M;
input  MMUART_1_RI_F2M;
input  MMUART_1_DSR_F2M;
input  MMUART_1_CTS_F2M;
input  MMUART_1_RXD_F2M;
input  MMUART_1_CLK_F2M;
input  MMUART_2_RXD_F2M;
input  MMUART_3_RXD_F2M;
input  MMUART_4_RXD_F2M;
input  CAN_0_RXBUS_F2M;
input  CAN_1_RXBUS_F2M;
input  CAN_CLK_F2M;
input  [3:0] QSPI_DATA_F2M;
input  SPI_0_SS_F2M;
input  SPI_0_DI_F2M;
input  SPI_0_CLK_F2M;
input  SPI_1_SS_F2M;
input  SPI_1_DI_F2M;
input  SPI_1_CLK_F2M;
input  I2C_0_SCL_F2M;
input  I2C_1_SCL_F2M;
input  I2C_0_SDA_F2M;
input  I2C_1_SDA_F2M;
input  I2C_0_BCLK_F2M;
input  I2C_0_SMBALERT_NI_F2M;
input  I2C_0_SMBSUS_NI_F2M;
input  I2C_1_BCLK_F2M;
input  I2C_1_SMBALERT_NI_F2M;
input  I2C_1_SMBSUS_NI_F2M;
input  [31:0] GPIO_2_F2M;
input  MAC_0_MDI_F2M;
input  MAC_1_MDI_F2M;
input  JTAG_TMS_F2M;
input  JTAG_TCK_F2M;
input  JTAG_TDI_F2M;
input  JTAG_TRSTB_F2M;
input  [63:0] MSS_INT_F2M;
input  [37:0] SPARE_1_F2M;
input  [37:0] SPARE_2_F2M;
input  BOOT_FAIL_CLEAR_F2M;
input  MSS_RESET_N_F2M;
input  GPIO_RESET_N_F2M;
input  USOC_TRACE_CLOCK_F2M;
input  USOC_TRACE_VALID_F2M;
input  [39:0] USOC_TRACE_DATA_F2M;
input  SPARE_5_F2M;
input  [7:0] MAC_0_GMII_MII_RXD_F2M;
input  MAC_0_GMII_MII_RX_DV_F2M;
input  MAC_0_GMII_MII_RX_ER_F2M;
input  MAC_0_GMII_MII_RX_CRS_F2M;
input  MAC_0_GMII_MII_RX_COL_F2M;
input  MAC_0_GMII_MII_RX_CLK_F2M;
input  MAC_0_GMII_MII_TX_CLK_F2M;
input  MAC_0_TSU_CLK_F2M;
input  [7:0] MAC_1_GMII_MII_RXD_F2M;
input  MAC_1_GMII_MII_RX_DV_F2M;
input  MAC_1_GMII_MII_RX_ER_F2M;
input  MAC_1_GMII_MII_RX_CRS_F2M;
input  MAC_1_GMII_MII_RX_COL_F2M;
input  MAC_1_GMII_MII_RX_CLK_F2M;
input  MAC_1_GMII_MII_TX_CLK_F2M;
input  MAC_1_TSU_CLK_F2M;
input  MAC_0_FILTER_MATCH1_F2M;
input  MAC_0_FILTER_MATCH2_F2M;
input  MAC_0_FILTER_MATCH3_F2M;
input  MAC_0_FILTER_MATCH4_F2M;
input  MAC_1_FILTER_MATCH1_F2M;
input  MAC_1_FILTER_MATCH2_F2M;
input  MAC_1_FILTER_MATCH3_F2M;
input  MAC_1_FILTER_MATCH4_F2M;
input  MAC_0_TSU_GEM_MS_F2M;
input  [1:0] MAC_0_TSU_GEM_INC_CTRL_F2M;
input  MAC_1_TSU_GEM_MS_F2M;
input  [1:0] MAC_1_TSU_GEM_INC_CTRL_F2M;
input  CRYPTO_HCLK;
input  CRYPTO_HRESETN;
input  CRYPTO_AHB_M_HREADY;
input  CRYPTO_AHB_M_HRESP;
input  [31:0] CRYPTO_AHB_M_HRDATA;
input  CRYPTO_AHB_S_HSEL;
input  [16:0] CRYPTO_AHB_S_HADDR;
input  [31:0] CRYPTO_AHB_S_HWDATA;
input  [1:0] CRYPTO_AHB_S_HSIZE;
input  [1:0] CRYPTO_AHB_S_HTRANS;
input  CRYPTO_AHB_S_HWRITE;
input  CRYPTO_AHB_S_HREADY;
input  CRYPTO_STALL_F2M;
input  CRYPTO_PURGE_F2M;
input  CRYPTO_GO_F2M;
input  CRYPTO_REQUEST_F2M;
input  CRYPTO_RELEASE_F2M;
input  CRYPTO_XENABLE_F2M;
input  [31:0] CRYPTO_XWDATA_F2M;
input  CRYPTO_XOUTACK_F2M;
input  CRYPTO_MESH_CLEAR_F2M;
input  EMMC_SD_CLK_F2M;
output FIC_0_DLL_LOCK_M2F;
output FIC_1_DLL_LOCK_M2F;
output FIC_2_DLL_LOCK_M2F;
output FIC_3_DLL_LOCK_M2F;
output [7:0] FIC_0_AXI4_M_AWID;
output [37:0] FIC_0_AXI4_M_AWADDR;
output [7:0] FIC_0_AXI4_M_AWLEN;
output [2:0] FIC_0_AXI4_M_AWSIZE;
output [1:0] FIC_0_AXI4_M_AWBURST;
output FIC_0_AXI4_M_AWLOCK;
output [3:0] FIC_0_AXI4_M_AWQOS;
output [3:0] FIC_0_AXI4_M_AWCACHE;
output [2:0] FIC_0_AXI4_M_AWPROT;
output FIC_0_AXI4_M_AWVALID;
output [63:0] FIC_0_AXI4_M_WDATA;
output [7:0] FIC_0_AXI4_M_WSTRB;
output FIC_0_AXI4_M_WLAST;
output FIC_0_AXI4_M_WVALID;
output FIC_0_AXI4_M_BREADY;
output [7:0] FIC_0_AXI4_M_ARID;
output [37:0] FIC_0_AXI4_M_ARADDR;
output [7:0] FIC_0_AXI4_M_ARLEN;
output [2:0] FIC_0_AXI4_M_ARSIZE;
output [1:0] FIC_0_AXI4_M_ARBURST;
output FIC_0_AXI4_M_ARLOCK;
output [3:0] FIC_0_AXI4_M_ARQOS;
output [3:0] FIC_0_AXI4_M_ARCACHE;
output [2:0] FIC_0_AXI4_M_ARPROT;
output FIC_0_AXI4_M_ARVALID;
output FIC_0_AXI4_M_RREADY;
output FIC_0_AXI4_S_AWREADY;
output FIC_0_AXI4_S_WREADY;
output [3:0] FIC_0_AXI4_S_BID;
output [1:0] FIC_0_AXI4_S_BRESP;
output FIC_0_AXI4_S_BVALID;
output FIC_0_AXI4_S_ARREADY;
output [3:0] FIC_0_AXI4_S_RID;
output [63:0] FIC_0_AXI4_S_RDATA;
output [1:0] FIC_0_AXI4_S_RRESP;
output FIC_0_AXI4_S_RLAST;
output FIC_0_AXI4_S_RVALID;
output [7:0] FIC_1_AXI4_M_AWID;
output [37:0] FIC_1_AXI4_M_AWADDR;
output [7:0] FIC_1_AXI4_M_AWLEN;
output [2:0] FIC_1_AXI4_M_AWSIZE;
output [1:0] FIC_1_AXI4_M_AWBURST;
output FIC_1_AXI4_M_AWLOCK;
output [3:0] FIC_1_AXI4_M_AWQOS;
output [3:0] FIC_1_AXI4_M_AWCACHE;
output [2:0] FIC_1_AXI4_M_AWPROT;
output FIC_1_AXI4_M_AWVALID;
output [63:0] FIC_1_AXI4_M_WDATA;
output [7:0] FIC_1_AXI4_M_WSTRB;
output FIC_1_AXI4_M_WLAST;
output FIC_1_AXI4_M_WVALID;
output FIC_1_AXI4_M_BREADY;
output [7:0] FIC_1_AXI4_M_ARID;
output [37:0] FIC_1_AXI4_M_ARADDR;
output [7:0] FIC_1_AXI4_M_ARLEN;
output [2:0] FIC_1_AXI4_M_ARSIZE;
output [1:0] FIC_1_AXI4_M_ARBURST;
output FIC_1_AXI4_M_ARLOCK;
output [3:0] FIC_1_AXI4_M_ARQOS;
output [3:0] FIC_1_AXI4_M_ARCACHE;
output [2:0] FIC_1_AXI4_M_ARPROT;
output FIC_1_AXI4_M_ARVALID;
output FIC_1_AXI4_M_RREADY;
output FIC_1_AXI4_S_AWREADY;
output FIC_1_AXI4_S_WREADY;
output [3:0] FIC_1_AXI4_S_BID;
output [1:0] FIC_1_AXI4_S_BRESP;
output FIC_1_AXI4_S_BVALID;
output FIC_1_AXI4_S_ARREADY;
output [3:0] FIC_1_AXI4_S_RID;
output [63:0] FIC_1_AXI4_S_RDATA;
output [1:0] FIC_1_AXI4_S_RRESP;
output FIC_1_AXI4_S_RLAST;
output FIC_1_AXI4_S_RVALID;
output FIC_2_AXI4_S_AWREADY;
output FIC_2_AXI4_S_WREADY;
output [3:0] FIC_2_AXI4_S_BID;
output [1:0] FIC_2_AXI4_S_BRESP;
output FIC_2_AXI4_S_BVALID;
output FIC_2_AXI4_S_ARREADY;
output [3:0] FIC_2_AXI4_S_RID;
output [63:0] FIC_2_AXI4_S_RDATA;
output [1:0] FIC_2_AXI4_S_RRESP;
output FIC_2_AXI4_S_RLAST;
output FIC_2_AXI4_S_RVALID;
output FIC_3_APB_M_PSEL;
output [28:0] FIC_3_APB_M_PADDR;
output FIC_3_APB_M_PWRITE;
output FIC_3_APB_M_PENABLE;
output [3:0] FIC_3_APB_M_PSTRB;
output [31:0] FIC_3_APB_M_PWDATA;
output MMUART_0_DTR_M2F;
output MMUART_0_RTS_M2F;
output MMUART_0_TXD_M2F;
output MMUART_0_TXD_OE_M2F;
output MMUART_1_DTR_M2F;
output MMUART_1_RTS_M2F;
output MMUART_1_TXD_M2F;
output MMUART_1_TXD_OE_M2F;
output MMUART_0_OUT1N_M2F;
output MMUART_0_OUT2N_M2F;
output MMUART_0_TE_M2F;
output MMUART_0_ESWM_M2F;
output MMUART_0_CLK_M2F;
output MMUART_0_CLK_OE_M2F;
output MMUART_1_OUT1N_M2F;
output MMUART_1_OUT2N_M2F;
output MMUART_1_TE_M2F;
output MMUART_1_ESWM_M2F;
output MMUART_1_CLK_M2F;
output MMUART_1_CLK_OE_M2F;
output MMUART_2_TXD_M2F;
output MMUART_3_TXD_M2F;
output MMUART_4_TXD_M2F;
output CAN_0_TX_EBL_M2F;
output CAN_0_TXBUS_M2F;
output CAN_1_TX_EBL_M2F;
output CAN_1_TXBUS_M2F;
output QSPI_SEL_M2F;
output QSPI_SEL_OE_M2F;
output QSPI_CLK_M2F;
output QSPI_CLK_OE_M2F;
output [3:0] QSPI_DATA_M2F;
output [3:0] QSPI_DATA_OE_M2F;
output SPI_0_SS1_M2F;
output SPI_0_SS1_OE_M2F;
output SPI_1_SS1_M2F;
output SPI_1_SS1_OE_M2F;
output SPI_0_DO_M2F;
output SPI_0_DO_OE_M2F;
output SPI_0_CLK_M2F;
output SPI_0_CLK_OE_M2F;
output SPI_1_DO_M2F;
output SPI_1_DO_OE_M2F;
output SPI_1_CLK_M2F;
output SPI_1_CLK_OE_M2F;
output I2C_0_SCL_OE_M2F;
output I2C_0_SDA_OE_M2F;
output I2C_1_SCL_OE_M2F;
output I2C_1_SDA_OE_M2F;
output I2C_0_SMBALERT_NO_M2F;
output I2C_0_SMBSUS_NO_M2F;
output I2C_1_SMBALERT_NO_M2F;
output I2C_1_SMBSUS_NO_M2F;
output [31:0] GPIO_2_M2F;
output [31:0] GPIO_2_OE_M2F;
output MAC_0_MDO_M2F;
output MAC_0_MDO_OE_M2F;
output MAC_0_MDC_M2F;
output MAC_1_MDO_M2F;
output MAC_1_MDO_OE_M2F;
output MAC_1_MDC_M2F;
output JTAG_TDO_M2F;
output JTAG_TDO_OE_M2F;
output [15:0] MSS_INT_M2F;
output [37:0] SPARE_M2F;
output PLL_CPU_LOCK_M2F;
output PLL_DDR_LOCK_M2F;
output PLL_SGMII_LOCK_M2F;
output [16:0] MSS_STATUS_M2F;
output BOOT_FAIL_ERROR_M2F;
output MSS_RESET_N_M2F;
output [4:0] SPARE_2_M2F;
output SPARE_3_M2F;
output [2:0] SPARE_4_M2F;
output [6:0] SPARE_5_M2F;
output WDOG_0_INTERRUPT_M2F;
output WDOG_1_INTERRUPT_M2F;
output WDOG_2_INTERRUPT_M2F;
output WDOG_3_INTERRUPT_M2F;
output WDOG_4_INTERRUPT_M2F;
output MPU_VIOLATION_FROM_FIC_0_M2F;
output MPU_VIOLATION_FROM_FIC_1_M2F;
output MPU_VIOLATION_FROM_FIC_2_M2F;
output MPU_VIOLATION_FROM_CRYPTO_M2F;
output MPU_VIOLATION_FROM_MAC_0_M2F;
output MPU_VIOLATION_FROM_MAC_1_M2F;
output MPU_VIOLATION_FROM_USB_M2F;
output MPU_VIOLATION_FROM_EMMC_SD_M2F;
output MPU_VIOLATION_FROM_SCB_M2F;
output MPU_VIOLATION_FROM_TRACE_M2F;
output REBOOT_REQUESTED_M2F;
output CPU_IN_RESET_M2F;
output AXI_IN_RESET_M2F;
output SCB_PERIPH_RESET_OCCURRED_M2F;
output SCB_MSS_RESET_OCCURRED_M2F;
output SCB_CPU_RESET_OCCURRED_M2F;
output DEBUGGER_RESET_OCCURRED_M2F;
output FABRIC_RESET_OCCURRED_M2F;
output WDOG_RESET_OCCURRED_M2F;
output GPIO_RESET_OCCURRED_M2F;
output SCB_BUS_RESET_OCCURRED_M2F;
output CPU_SOFT_RESET_OCCURRED_M2F;
output [1:0] CPU_CLK_DIVIDER_M2F;
output [1:0] AXI_CLK_DIVIDER_M2F;
output [1:0] AHB_APB_CLK_DIVIDER_M2F;
output [7:0] USOC_CONTROL_DATA_M2F;
output [7:0] MAC_0_GMII_MII_TXD_M2F;
output MAC_0_GMII_MII_TX_EN_M2F;
output MAC_0_GMII_MII_TX_ER_M2F;
output MAC_0_LOCAL_LOOPBACK_M2F;
output MAC_0_LOOPBACK_M2F;
output MAC_0_HALF_DUPLEX_M2F;
output [3:0] MAC_0_SPEED_MODE_M2F;
output [7:0] MAC_1_GMII_MII_TXD_M2F;
output MAC_1_GMII_MII_TX_EN_M2F;
output MAC_1_GMII_MII_TX_ER_M2F;
output MAC_1_LOCAL_LOOPBACK_M2F;
output MAC_1_LOOPBACK_M2F;
output MAC_1_HALF_DUPLEX_M2F;
output [3:0] MAC_1_SPEED_MODE_M2F;
output [127:0] MAC_0_FILTER_DATA_M2F;
output MAC_0_FILTER_SA_STB_M2F;
output MAC_0_FILTER_DA_STB_M2F;
output MAC_0_FILTER_TYPE_STB_M2F;
output MAC_0_FILTER_VLAN_TAG1_STB_M2F;
output MAC_0_FILTER_VLAN_TAG2_STB_M2F;
output MAC_0_FILTER_IP_SA_STB_M2F;
output MAC_0_FILTER_IP_DA_STB_M2F;
output MAC_0_FILTER_SP_STB_M2F;
output MAC_0_FILTER_DP_STB_M2F;
output MAC_0_FILTER_IPV6_M2F;
output MAC_0_WOL_M2F;
output [127:0] MAC_1_FILTER_DATA_M2F;
output MAC_1_FILTER_SA_STB_M2F;
output MAC_1_FILTER_DA_STB_M2F;
output MAC_1_FILTER_TYPE_STB_M2F;
output MAC_1_FILTER_VLAN_TAG1_STB_M2F;
output MAC_1_FILTER_VLAN_TAG2_STB_M2F;
output MAC_1_FILTER_IP_SA_STB_M2F;
output MAC_1_FILTER_IP_DA_STB_M2F;
output MAC_1_FILTER_SP_STB_M2F;
output MAC_1_FILTER_DP_STB_M2F;
output MAC_1_FILTER_IPV6_M2F;
output MAC_1_WOL_M2F;
output MAC_0_TSU_SOF_TX_M2F;
output MAC_0_TSU_SYNC_FRAME_TX_M2F;
output MAC_0_TSU_DELAY_REQ_TX_M2F;
output MAC_0_TSU_PDELAY_REQ_TX_M2F;
output MAC_0_TSU_PDELAY_RESP_TX_M2F;
output MAC_0_TSU_SOF_RX_M2F;
output MAC_0_TSU_SYNC_FRAME_RX_M2F;
output MAC_0_TSU_DELAY_REQ_RX_M2F;
output MAC_0_TSU_PDELAY_REQ_RX_M2F;
output MAC_0_TSU_PDELAY_RESP_RX_M2F;
output [93:0] MAC_0_TSU_TIMER_CNT_M2F;
output MAC_0_TSU_TIMER_CMP_VAL_M2F;
output MAC_1_TSU_SOF_TX_M2F;
output MAC_1_TSU_SYNC_FRAME_TX_M2F;
output MAC_1_TSU_DELAY_REQ_TX_M2F;
output MAC_1_TSU_PDELAY_REQ_TX_M2F;
output MAC_1_TSU_PDELAY_RESP_TX_M2F;
output MAC_1_TSU_SOF_RX_M2F;
output MAC_1_TSU_SYNC_FRAME_RX_M2F;
output MAC_1_TSU_DELAY_REQ_RX_M2F;
output MAC_1_TSU_PDELAY_REQ_RX_M2F;
output MAC_1_TSU_PDELAY_RESP_RX_M2F;
output [93:0] MAC_1_TSU_TIMER_CNT_M2F;
output MAC_1_TSU_TIMER_CMP_VAL_M2F;
output CRYPTO_DLL_LOCK_M2F;
output [31:0] CRYPTO_AHB_M_HADDR;
output [31:0] CRYPTO_AHB_M_HWDATA;
output [1:0] CRYPTO_AHB_M_HSIZE;
output [1:0] CRYPTO_AHB_M_HTRANS;
output CRYPTO_AHB_M_HWRITE;
output CRYPTO_AHB_M_HMASTLOCK;
output CRYPTO_AHB_S_HREADYOUT;
output CRYPTO_AHB_S_HRESP;
output [31:0] CRYPTO_AHB_S_HRDATA;
output CRYPTO_BUSY_M2F;
output CRYPTO_COMPLETE_M2F;
output CRYPTO_ALARM_M2F;
output CRYPTO_BUSERROR_M2F;
output CRYPTO_MSS_REQUEST_M2F;
output CRYPTO_MSS_RELEASE_M2F;
output CRYPTO_OWNER_M2F;
output CRYPTO_MSS_OWNER_M2F;
output [9:0] CRYPTO_XWADDR_M2F;
output CRYPTO_XINACCEPT_M2F;
output [31:0] CRYPTO_XRDATA_M2F;
output [9:0] CRYPTO_XRADDR_M2F;
output CRYPTO_XVALIDOUT_M2F;
output CRYPTO_MESH_ERROR_M2F;
input  MSSIO37_IN;
output MSSIO37_OUT;
output MSSIO37_OE;
input  MSSIO36_IN;
output MSSIO36_OUT;
output MSSIO36_OE;
input  MSSIO35_IN;
output MSSIO35_OUT;
output MSSIO35_OE;
input  MSSIO34_IN;
output MSSIO34_OUT;
output MSSIO34_OE;
input  MSSIO33_IN;
output MSSIO33_OUT;
output MSSIO33_OE;
input  MSSIO32_IN;
output MSSIO32_OUT;
output MSSIO32_OE;
input  MSSIO31_IN;
output MSSIO31_OUT;
output MSSIO31_OE;
input  MSSIO30_IN;
output MSSIO30_OUT;
output MSSIO30_OE;
input  MSSIO29_IN;
output MSSIO29_OUT;
output MSSIO29_OE;
input  MSSIO28_IN;
output MSSIO28_OUT;
output MSSIO28_OE;
input  MSSIO27_IN;
output MSSIO27_OUT;
output MSSIO27_OE;
input  MSSIO26_IN;
output MSSIO26_OUT;
output MSSIO26_OE;
input  MSSIO25_IN;
output MSSIO25_OUT;
output MSSIO25_OE;
input  MSSIO24_IN;
output MSSIO24_OUT;
output MSSIO24_OE;
input  MSSIO23_IN;
output MSSIO23_OUT;
output MSSIO23_OE;
input  MSSIO22_IN;
output MSSIO22_OUT;
output MSSIO22_OE;
input  MSSIO21_IN;
output MSSIO21_OUT;
output MSSIO21_OE;
input  MSSIO20_IN;
output MSSIO20_OUT;
output MSSIO20_OE;
input  MSSIO19_IN;
output MSSIO19_OUT;
output MSSIO19_OE;
input  MSSIO18_IN;
output MSSIO18_OUT;
output MSSIO18_OE;
input  MSSIO17_IN;
output MSSIO17_OUT;
output MSSIO17_OE;
input  MSSIO16_IN;
output MSSIO16_OUT;
output MSSIO16_OE;
input  MSSIO15_IN;
output MSSIO15_OUT;
output MSSIO15_OE;
input  MSSIO14_IN;
output MSSIO14_OUT;
output MSSIO14_OE;
input  MSSIO13_IN;
output MSSIO13_OUT;
output MSSIO13_OE;
input  MSSIO12_IN;
output MSSIO12_OUT;
output MSSIO12_OE;
input  MSSIO11_IN;
output MSSIO11_OUT;
output MSSIO11_OE;
input  MSSIO10_IN;
output MSSIO10_OUT;
output MSSIO10_OE;
input  MSSIO9_IN;
output MSSIO9_OUT;
output MSSIO9_OE;
input  MSSIO8_IN;
output MSSIO8_OUT;
output MSSIO8_OE;
input  MSSIO7_IN;
output MSSIO7_OUT;
output MSSIO7_OE;
input  MSSIO6_IN;
output MSSIO6_OUT;
output MSSIO6_OE;
input  MSSIO5_IN;
output MSSIO5_OUT;
output MSSIO5_OE;
input  MSSIO4_IN;
output MSSIO4_OUT;
output MSSIO4_OE;
input  MSSIO3_IN;
output MSSIO3_OUT;
output MSSIO3_OE;
input  MSSIO2_IN;
output MSSIO2_OUT;
output MSSIO2_OE;
input  MSSIO1_IN;
output MSSIO1_OUT;
output MSSIO1_OE;
input  MSSIO0_IN;
output MSSIO0_OUT;
output MSSIO0_OE;
input  REFCLK;
input  SGMII_RX1;
input  SGMII_RX0;
output SGMII_TX1;
output SGMII_TX0;
input  DDR_DQS4_IN;
output DDR_DQS4_OUT;
output DDR_DQS4_OE;
input  DDR_DQS3_IN;
output DDR_DQS3_OUT;
output DDR_DQS3_OE;
input  DDR_DQS2_IN;
output DDR_DQS2_OUT;
output DDR_DQS2_OE;
input  DDR_DQS1_IN;
output DDR_DQS1_OUT;
output DDR_DQS1_OE;
input  DDR_DQS0_IN;
output DDR_DQS0_OUT;
output DDR_DQS0_OE;
output DDR_CK1;
output DDR_CK0;
output DDR3_WE_N;
output DDR_PARITY;
output DDR_RAM_RST_N;
input  DDR_ALERT_N;
output DDR_ACT_N;
output DDR_A16;
output DDR_A15;
output DDR_A14;
output DDR_A13;
output DDR_A12;
output DDR_A11;
output DDR_A10;
output DDR_A9;
output DDR_A8;
output DDR_A7;
output DDR_A6;
output DDR_A5;
output DDR_A4;
output DDR_A3;
output DDR_A2;
output DDR_A1;
output DDR_A0;
output DDR_BA1;
output DDR_BA0;
output DDR_BG1;
output DDR_BG0;
output DDR_CKE1;
output DDR_CKE0;
output DDR_CS1;
output DDR_CS0;
output DDR_ODT1;
output DDR_ODT0;
input  DDR_DQ35_IN;
output DDR_DQ35_OUT;
output DDR_DQ35_OE;
input  DDR_DQ34_IN;
output DDR_DQ34_OUT;
output DDR_DQ34_OE;
input  DDR_DQ33_IN;
output DDR_DQ33_OUT;
output DDR_DQ33_OE;
input  DDR_DQ32_IN;
output DDR_DQ32_OUT;
output DDR_DQ32_OE;
input  DDR_DQ31_IN;
output DDR_DQ31_OUT;
output DDR_DQ31_OE;
input  DDR_DQ30_IN;
output DDR_DQ30_OUT;
output DDR_DQ30_OE;
input  DDR_DQ29_IN;
output DDR_DQ29_OUT;
output DDR_DQ29_OE;
input  DDR_DQ28_IN;
output DDR_DQ28_OUT;
output DDR_DQ28_OE;
input  DDR_DQ27_IN;
output DDR_DQ27_OUT;
output DDR_DQ27_OE;
input  DDR_DQ26_IN;
output DDR_DQ26_OUT;
output DDR_DQ26_OE;
input  DDR_DQ25_IN;
output DDR_DQ25_OUT;
output DDR_DQ25_OE;
input  DDR_DQ24_IN;
output DDR_DQ24_OUT;
output DDR_DQ24_OE;
input  DDR_DQ23_IN;
output DDR_DQ23_OUT;
output DDR_DQ23_OE;
input  DDR_DQ22_IN;
output DDR_DQ22_OUT;
output DDR_DQ22_OE;
input  DDR_DQ21_IN;
output DDR_DQ21_OUT;
output DDR_DQ21_OE;
input  DDR_DQ20_IN;
output DDR_DQ20_OUT;
output DDR_DQ20_OE;
input  DDR_DQ19_IN;
output DDR_DQ19_OUT;
output DDR_DQ19_OE;
input  DDR_DQ18_IN;
output DDR_DQ18_OUT;
output DDR_DQ18_OE;
input  DDR_DQ17_IN;
output DDR_DQ17_OUT;
output DDR_DQ17_OE;
input  DDR_DQ16_IN;
output DDR_DQ16_OUT;
output DDR_DQ16_OE;
input  DDR_DQ15_IN;
output DDR_DQ15_OUT;
output DDR_DQ15_OE;
input  DDR_DQ14_IN;
output DDR_DQ14_OUT;
output DDR_DQ14_OE;
input  DDR_DQ13_IN;
output DDR_DQ13_OUT;
output DDR_DQ13_OE;
input  DDR_DQ12_IN;
output DDR_DQ12_OUT;
output DDR_DQ12_OE;
input  DDR_DQ11_IN;
output DDR_DQ11_OUT;
output DDR_DQ11_OE;
input  DDR_DQ10_IN;
output DDR_DQ10_OUT;
output DDR_DQ10_OE;
input  DDR_DQ9_IN;
output DDR_DQ9_OUT;
output DDR_DQ9_OE;
input  DDR_DQ8_IN;
output DDR_DQ8_OUT;
output DDR_DQ8_OE;
input  DDR_DQ7_IN;
output DDR_DQ7_OUT;
output DDR_DQ7_OE;
input  DDR_DQ6_IN;
output DDR_DQ6_OUT;
output DDR_DQ6_OE;
input  DDR_DQ5_IN;
output DDR_DQ5_OUT;
output DDR_DQ5_OE;
input  DDR_DQ4_IN;
output DDR_DQ4_OUT;
output DDR_DQ4_OE;
input  DDR_DQ3_IN;
output DDR_DQ3_OUT;
output DDR_DQ3_OE;
input  DDR_DQ2_IN;
output DDR_DQ2_OUT;
output DDR_DQ2_OE;
input  DDR_DQ1_IN;
output DDR_DQ1_OUT;
output DDR_DQ1_OE;
input  DDR_DQ0_IN;
output DDR_DQ0_OUT;
output DDR_DQ0_OE;
input  DDR_DM0_IN;
output DDR_DM0_OUT;
output DDR_DM0_OE;
input  DDR_DM1_IN;
output DDR_DM1_OUT;
output DDR_DM1_OE;
input  DDR_DM2_IN;
output DDR_DM2_OUT;
output DDR_DM2_OE;
input  DDR_DM3_IN;
output DDR_DM3_OUT;
output DDR_DM3_OE;
input  DDR_DM4_IN;
output DDR_DM4_OUT;
output DDR_DM4_OE;
input  REFCLK_0_PLL_NW;
input  REFCLK_1_PLL_NW;
parameter CRYPTO_MODE = "";
parameter BOOT_MODE = "";
parameter BOOT_MODE1_E51_START_ADDRESS_ENVM = 'h0;
parameter BOOT_MODE1_U54_1_START_ADDRESS_ENVM = 'h0;
parameter BOOT_MODE1_U54_2_START_ADDRESS_ENVM = 'h0;
parameter BOOT_MODE1_U54_3_START_ADDRESS_ENVM = 'h0;
parameter BOOT_MODE1_U54_4_START_ADDRESS_ENVM = 'h0;
parameter BOOT_MODE2_START_PAGE_SNVM = 0;
parameter BOOT_MODE3_START_ADDRESS_ENVM = 'h0;
parameter MSS_CLK_DIV = 0;
parameter MSS_AHB_APB_CLK_DIV = 0;
parameter MSS_AXI_CLK_DIV = 0;
parameter MSS_CLK_FREQ = 0.0;
parameter CRYPTO_MSS_CLK_FREQ = 0.0;
parameter MSS_DDR_CLK_FREQ = 0.0;
parameter PROGRAM_NAME = "";
parameter CORE_NAME = "";
parameter DIE = "";
parameter PKG = "";
parameter BANK2_VDDI = "";
parameter BANK4_VDDI = "";
parameter BANK5_VDDI = "";
parameter DDR_SDRAM_TYPE = "";
parameter REFCLK_IOSTD = "";
parameter SGMII_IOSTD = "";
parameter SGMII_RX0_IOSTD = "";
parameter SGMII_RX1_IOSTD = "";
parameter SGMII_TX0_IOSTD = "";
parameter SGMII_TX1_IOSTD = "";
parameter SPI0_CONTROL1_CFG_MODE = 'h0;
parameter SPI1_CONTROL1_CFG_MODE = 'h0;
parameter DDR_SEGS_SEG0_0_ADDRESS_OFFSET = 'h7F80;
parameter DDR_SEGS_SEG0_1_ADDRESS_OFFSET = 'h7000;
parameter DDR_SEGS_SEG1_2_ADDRESS_OFFSET = 'h7F40;
parameter DDR_SEGS_SEG1_3_ADDRESS_OFFSET = 'h6C00;
parameter DDR_SEGS_SEG1_4_ADDRESS_OFFSET = 'h7F30;
parameter DDR_SEGS_SEG1_5_ADDRESS_OFFSET = 'h6800;
parameter DDR_SEGS_SEG1_6_ADDRESS_OFFSET = 'h0;
parameter DDR_DDRC_CFG_AXI_START_ADDRESS_AXI1_0 = 'h0;
parameter DDR_DDRC_CFG_AXI_START_ADDRESS_AXI1_1 = 'h0;
parameter DDR_DDRC_CFG_AXI_START_ADDRESS_AXI2_0 = 'h0;
parameter DDR_DDRC_CFG_AXI_START_ADDRESS_AXI2_1 = 'h0;
parameter DDR_DDRC_CFG_AXI_END_ADDRESS_AXI1_0 = 'hFFFFFFFF;
parameter DDR_DDRC_CFG_AXI_END_ADDRESS_AXI1_1 = 'h3;
parameter DDR_DDRC_CFG_AXI_END_ADDRESS_AXI2_0 = 'hFFFFFFFF;
parameter DDR_DDRC_CFG_AXI_END_ADDRESS_AXI2_1 = 'h3;
parameter DDR_DDRC_CFG_MEM_START_ADDRESS_AXI1_0 = 'h0;
parameter DDR_DDRC_CFG_MEM_START_ADDRESS_AXI1_1 = 'h0;
parameter DDR_DDRC_CFG_MEM_START_ADDRESS_AXI2_0 = 'h0;
parameter DDR_DDRC_CFG_MEM_START_ADDRESS_AXI2_1 = 'h0;
parameter MSSIO_IOMUX0_CR_SPI0_FABRIC = 'h0;
parameter MSSIO_IOMUX0_CR_SPI1_FABRIC = 'h0;
parameter MSSIO_IOMUX0_CR_I2C0_FABRIC = 'h0;
parameter MSSIO_IOMUX0_CR_I2C1_FABRIC = 'h0;
parameter MSSIO_IOMUX0_CR_CAN0_FABRIC = 'h0;
parameter MSSIO_IOMUX0_CR_CAN1_FABRIC = 'h0;
parameter MSSIO_IOMUX0_CR_QSPI_FABRIC = 'h0;
parameter MSSIO_IOMUX0_CR_MMUART0_FABRIC = 'h0;
parameter MSSIO_IOMUX0_CR_MMUART1_FABRIC = 'h0;
parameter MSSIO_IOMUX0_CR_MMUART2_FABRIC = 'h0;
parameter MSSIO_IOMUX0_CR_MMUART3_FABRIC = 'h0;
parameter MSSIO_IOMUX0_CR_MMUART4_FABRIC = 'h0;
parameter MSSIO_IOMUX0_CR_MDIO0_FABRIC = 'h0;
parameter MSSIO_IOMUX0_CR_MDIO1_FABRIC = 'h0;
parameter MSSIO_IOMUX1_CR_PAD0 = 'hF;
parameter MSSIO_IOMUX1_CR_PAD1 = 'hF;
parameter MSSIO_IOMUX1_CR_PAD2 = 'hF;
parameter MSSIO_IOMUX1_CR_PAD3 = 'hF;
parameter MSSIO_IOMUX1_CR_PAD4 = 'hF;
parameter MSSIO_IOMUX1_CR_PAD5 = 'hF;
parameter MSSIO_IOMUX1_CR_PAD6 = 'hF;
parameter MSSIO_IOMUX1_CR_PAD7 = 'hF;
parameter MSSIO_IOMUX2_CR_PAD8 = 'hF;
parameter MSSIO_IOMUX2_CR_PAD9 = 'hF;
parameter MSSIO_IOMUX2_CR_PAD10 = 'hF;
parameter MSSIO_IOMUX2_CR_PAD11 = 'hF;
parameter MSSIO_IOMUX2_CR_PAD12 = 'hF;
parameter MSSIO_IOMUX2_CR_PAD13 = 'hF;
parameter MSSIO_IOMUX3_CR_PAD14 = 'hF;
parameter MSSIO_IOMUX3_CR_PAD15 = 'hF;
parameter MSSIO_IOMUX3_CR_PAD16 = 'hF;
parameter MSSIO_IOMUX3_CR_PAD17 = 'hF;
parameter MSSIO_IOMUX3_CR_PAD18 = 'hF;
parameter MSSIO_IOMUX3_CR_PAD19 = 'hF;
parameter MSSIO_IOMUX3_CR_PAD20 = 'hF;
parameter MSSIO_IOMUX3_CR_PAD21 = 'hF;
parameter MSSIO_IOMUX4_CR_PAD22 = 'hF;
parameter MSSIO_IOMUX4_CR_PAD23 = 'hF;
parameter MSSIO_IOMUX4_CR_PAD24 = 'hF;
parameter MSSIO_IOMUX4_CR_PAD25 = 'hF;
parameter MSSIO_IOMUX4_CR_PAD26 = 'hF;
parameter MSSIO_IOMUX4_CR_PAD27 = 'hF;
parameter MSSIO_IOMUX4_CR_PAD28 = 'hF;
parameter MSSIO_IOMUX4_CR_PAD29 = 'hF;
parameter MSSIO_IOMUX5_CR_PAD30 = 'hF;
parameter MSSIO_IOMUX5_CR_PAD31 = 'hF;
parameter MSSIO_IOMUX5_CR_PAD32 = 'hF;
parameter MSSIO_IOMUX5_CR_PAD33 = 'hF;
parameter MSSIO_IOMUX5_CR_PAD34 = 'hF;
parameter MSSIO_IOMUX5_CR_PAD35 = 'hF;
parameter MSSIO_IOMUX5_CR_PAD36 = 'hF;
parameter MSSIO_IOMUX5_CR_PAD37 = 'hF;
parameter MSSIO_IOMUX6_CR_VLT_SEL = 'h0;
parameter MSSIO_IOMUX6_CR_VLT_EN = 'h0;
parameter MSSIO_IOMUX6_CR_VLT_CMD_DIR = 'h0;
parameter MSSIO_IOMUX6_CR_VLT_DIR_0 = 'h0;
parameter MSSIO_IOMUX6_CR_VLT_DIR_1_3 = 'h0;
parameter MSSIO_IOMUX6_CR_SD_LED = 'h0;
parameter MSSIO_IOMUX6_CR_SD_VOLT_0 = 'h0;
parameter MSSIO_IOMUX6_CR_SD_VOLT_1 = 'h0;
parameter MSSIO_IOMUX6_CR_SD_VOLT_2 = 'h0;
parameter MSSIO_MSSIO_BANK2_CFG_CR_BANK_PCODE = 'h7;
parameter MSSIO_MSSIO_BANK2_CFG_CR_BANK_NCODE = 'h9;
parameter MSSIO_MSSIO_BANK2_CFG_CR_VS = 'h8;
parameter MSSIO_MSSIO_BANK4_CFG_CR_BANK_PCODE = 'h7;
parameter MSSIO_MSSIO_BANK4_CFG_CR_BANK_NCODE = 'h9;
parameter MSSIO_MSSIO_BANK4_CFG_CR_VS = 'h8;
parameter SGMII_SGMII_MODE_REG_BC_VS = 'h8;
parameter SGMII_SGMII_MODE_REG_PLL_EN = 'h0;
parameter SGMII_SGMII_MODE_REG_DLL_EN = 'h0;
parameter SGMII_DYN_CNTL_REG_PLL_SOFT_RESET_PERIPH = 'h0;
parameter SGMII_DYN_CNTL_REG_DLL_SOFT_RESET_PERIPH = 'h0;
parameter SGMII_DYN_CNTL_REG_PVT_SOFT_RESET_PERIPH = 'h1;
parameter SGMII_DYN_CNTL_REG_BC_SOFT_RESET_PERIPH = 'h0;
parameter SGMII_SGMII_MODE_REG_TX0_EN = 'h0;
parameter SGMII_SGMII_MODE_REG_RX0_EN = 'h0;
parameter SGMII_SGMII_MODE_REG_CH0_CDR_RESET_B = 'h1;
parameter SGMII_DYN_CNTL_REG_LANE0_SOFT_RESET_PERIPH = 'h0;
parameter SGMII_CH0_CNTL_REG_TX0_WPU_P = 'h0;
parameter SGMII_CH0_CNTL_REG_TX0_WPD_P = 'h0;
parameter SGMII_CH0_CNTL_REG_TX0_SLEW_P = 'h0;
parameter SGMII_CH0_CNTL_REG_TX0_DRV_P = 'h0;
parameter SGMII_CH0_CNTL_REG_TX0_ODT_P = 'h0;
parameter SGMII_CH0_CNTL_REG_TX0_ODT_STATIC_P = 'h0;
parameter SGMII_CH0_CNTL_REG_RX0_WPU_P = 'h0;
parameter SGMII_CH0_CNTL_REG_RX0_WPD_P = 'h0;
parameter SGMII_CH0_CNTL_REG_RX0_IBUFMD_P = 'h7;
parameter SGMII_CH0_CNTL_REG_RX0_ODT_P = 'h0;
parameter SGMII_CH0_CNTL_REG_RX0_ODT_STATIC_P = 'h0;
parameter SGMII_SGMII_MODE_REG_TX1_EN = 'h0;
parameter SGMII_SGMII_MODE_REG_RX1_EN = 'h0;
parameter SGMII_SGMII_MODE_REG_CH1_CDR_RESET_B = 'h1;
parameter SGMII_DYN_CNTL_REG_LANE1_SOFT_RESET_PERIPH = 'h0;
parameter SGMII_CH1_CNTL_REG_TX1_WPU_P = 'h0;
parameter SGMII_CH1_CNTL_REG_TX1_WPD_P = 'h0;
parameter SGMII_CH1_CNTL_REG_TX1_SLEW_P = 'h0;
parameter SGMII_CH1_CNTL_REG_TX1_DRV_P = 'h0;
parameter SGMII_CH1_CNTL_REG_TX1_ODT_P = 'h0;
parameter SGMII_CH1_CNTL_REG_TX1_ODT_STATIC_P = 'h0;
parameter SGMII_CH1_CNTL_REG_RX1_WPU_P = 'h0;
parameter SGMII_CH1_CNTL_REG_RX1_WPD_P = 'h0;
parameter SGMII_CH1_CNTL_REG_RX1_IBUFMD_P = 'h7;
parameter SGMII_CH1_CNTL_REG_RX1_ODT_P = 'h0;
parameter SGMII_CH1_CNTL_REG_RX1_ODT_STATIC_P = 'h0;
parameter SGMII_SGMII_MODE_REG_PVT_EN = 'h1;
parameter SGMII_SGMII_MODE_REG_BC_VRGEN_EN = 'h1;
parameter SGMII_RECAL_CNTL_REG_PVT_CALIB_START = 'h1;
parameter SGMII_RECAL_CNTL_REG_PVT_CALIB_LOCK = 'h1;
parameter SGMII_DYN_CNTL_REG_CLKMUX_SOFT_RESET_PERIPH = 'h0;
parameter SGMII_CLK_CNTL_REG_REFCLK_EN_RXMODE_P = 'h3;
parameter SGMII_CLK_CNTL_REG_REFCLK_EN_RXMODE_N = 'h3;
parameter CLK_SGMII_CFM_CLK_XCVR_EN_RXMODE_P = 'h3;
parameter CLK_SGMII_CFM_CLK_XCVR_EN_RXMODE_N = 'h3;
parameter SGMII_SGMII_MODE_REG_REFCLK_EN_UDRIVE_P = 'h0;
parameter SGMII_SGMII_MODE_REG_REFCLK_EN_UDRIVE_N = 'h0;
parameter CLK_SGMII_CFM_CLK_XCVR_EN_UDRIVE_P = 'h0;
parameter CLK_SGMII_CFM_CLK_XCVR_EN_UDRIVE_N = 'h0;
parameter SGMII_SGMII_MODE_REG_REFCLK_EN_RDIFF = 'h1;
parameter CLK_SGMII_CFM_CLK_XCVR_EN_RDIFF = 'h1;
parameter SGMII_CLK_CNTL_REG_REFCLK_EN_TERM_P = 'h0;
parameter SGMII_CLK_CNTL_REG_REFCLK_EN_TERM_N = 'h0;
parameter CLK_SGMII_CFM_CLK_XCVR_EN_TERM_P = 'h0;
parameter CLK_SGMII_CFM_CLK_XCVR_EN_TERM_N = 'h0;
parameter SGMII_SGMII_MODE_REG_REFCLK_EN_INS_HYST_P = 'h0;
parameter SGMII_SGMII_MODE_REG_REFCLK_EN_INS_HYST_N = 'h0;
parameter CLK_SGMII_CFM_CLK_XCVR_EN_INS_HYST_P = 'h0;
parameter CLK_SGMII_CFM_CLK_XCVR_EN_INS_HYST_N = 'h0;
parameter SGMII_CLK_CNTL_REG_REFCLK_CLKBUF_EN_PULLUP = 'h0;
parameter CLK_SGMII_CFM_CLK_XCVR_CLKBUF_EN_PULLUP = 'h0;
parameter MSSIO_MSSIO_BANK4_IO_CFG_0_1_CR_IO_CFG_0 = 'h829;
parameter MSSIO_MSSIO_BANK4_IO_CFG_0_1_CR_IO_CFG_1 = 'h829;
parameter MSSIO_MSSIO_BANK4_IO_CFG_2_3_CR_IO_CFG_2 = 'h829;
parameter MSSIO_MSSIO_BANK4_IO_CFG_2_3_CR_IO_CFG_3 = 'h829;
parameter MSSIO_MSSIO_BANK4_IO_CFG_4_5_CR_IO_CFG_4 = 'h829;
parameter MSSIO_MSSIO_BANK4_IO_CFG_4_5_CR_IO_CFG_5 = 'h829;
parameter MSSIO_MSSIO_BANK4_IO_CFG_6_7_CR_IO_CFG_6 = 'h829;
parameter MSSIO_MSSIO_BANK4_IO_CFG_6_7_CR_IO_CFG_7 = 'h829;
parameter MSSIO_MSSIO_BANK4_IO_CFG_8_9_CR_IO_CFG_8 = 'h829;
parameter MSSIO_MSSIO_BANK4_IO_CFG_8_9_CR_IO_CFG_9 = 'h829;
parameter MSSIO_MSSIO_BANK4_IO_CFG_10_11_CR_IO_CFG_10 = 'h829;
parameter MSSIO_MSSIO_BANK4_IO_CFG_10_11_CR_IO_CFG_11 = 'h829;
parameter MSSIO_MSSIO_BANK4_IO_CFG_12_13_CR_IO_CFG_12 = 'h829;
parameter MSSIO_MSSIO_BANK4_IO_CFG_12_13_CR_IO_CFG_13 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_0_1_CR_IO_CFG_0 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_0_1_CR_IO_CFG_1 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_2_3_CR_IO_CFG_2 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_2_3_CR_IO_CFG_3 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_4_5_CR_IO_CFG_4 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_4_5_CR_IO_CFG_5 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_6_7_CR_IO_CFG_6 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_6_7_CR_IO_CFG_7 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_8_9_CR_IO_CFG_8 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_8_9_CR_IO_CFG_9 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_10_11_CR_IO_CFG_10 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_10_11_CR_IO_CFG_11 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_12_13_CR_IO_CFG_12 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_12_13_CR_IO_CFG_13 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_14_15_CR_IO_CFG_14 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_14_15_CR_IO_CFG_15 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_16_17_CR_IO_CFG_16 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_16_17_CR_IO_CFG_17 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_18_19_CR_IO_CFG_18 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_18_19_CR_IO_CFG_19 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_20_21_CR_IO_CFG_20 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_20_21_CR_IO_CFG_21 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_22_23_CR_IO_CFG_22 = 'h829;
parameter MSSIO_MSSIO_BANK2_IO_CFG_22_23_CR_IO_CFG_23 = 'h829;
parameter GENERAL_GPIO_CR_GPIO0_SOFT_RESET_SELECT = 'h3;
parameter GENERAL_GPIO_CR_GPIO1_SOFT_RESET_SELECT = 'h7;
parameter GENERAL_GPIO_CR_GPIO2_SOFT_RESET_SELECT = 'hF;
parameter GENERAL_CRYPTO_CR_INFO_MSS_MODE = 'h0;
parameter DDR_DDRC_CFG_CHIPADDR_MAP_CFG_CHIPADDR_MAP = 'h0;
parameter DDR_DDRC_CFG_BANKADDR_MAP_0_CFG_BANKADDR_MAP_0 = 'h0;
parameter DDR_DDRC_CFG_ROWADDR_MAP_0_CFG_ROWADDR_MAP_0 = 'h0;
parameter DDR_DDRC_CFG_ROWADDR_MAP_1_CFG_ROWADDR_MAP_1 = 'h0;
parameter DDR_DDRC_CFG_ROWADDR_MAP_2_CFG_ROWADDR_MAP_2 = 'h0;
parameter DDR_DDRC_CFG_ROWADDR_MAP_3_CFG_ROWADDR_MAP_3 = 'h0;
parameter DDR_DDRC_CFG_COLADDR_MAP_0_CFG_COLADDR_MAP_0 = 'h0;
parameter DDR_DDRC_CFG_COLADDR_MAP_1_CFG_COLADDR_MAP_1 = 'h0;
parameter DDR_DDRC_CFG_COLADDR_MAP_2_CFG_COLADDR_MAP_2 = 'h0;
parameter DDR_DDRC_CFG_MEM_COLBITS_CFG_MEM_COLBITS = 'hA;
parameter DDR_DDRC_CFG_MEM_ROWBITS_CFG_MEM_ROWBITS = 'hE;
parameter DDR_DDRC_CFG_MEM_BANKBITS_CFG_MEM_BANKBITS = 'h3;
parameter DDR_DDRC_CFG_CL_CFG_CL = 'hC;
parameter DDR_DDRC_CFG_CWL_CFG_CWL = 'hA;
parameter DDR_DDRC_CFG_NUM_RANKS_CFG_NUM_RANKS = 'h2;
parameter DDR_DDRC_CFG_ZQINIT_CAL_DURATION_CFG_ZQINIT_CAL_DURATION = 'h2AB;
parameter DDR_DDRC_CFG_ZQ_CAL_L_DURATION_CFG_ZQ_CAL_L_DURATION = 'h156;
parameter DDR_DDRC_CFG_ZQ_CAL_S_DURATION_CFG_ZQ_CAL_S_DURATION = 'h56;
parameter DDR_DDRC_CFG_ODT_RD_MAP_CS0_CFG_ODT_RD_MAP_CS0 = 'h2;
parameter DDR_DDRC_CFG_ODT_RD_MAP_CS1_CFG_ODT_RD_MAP_CS1 = 'h1;
parameter DDR_DDRC_CFG_ODT_WR_MAP_CS0_CFG_ODT_WR_MAP_CS0 = 'h1;
parameter DDR_DDRC_CFG_ODT_WR_MAP_CS1_CFG_ODT_WR_MAP_CS1 = 'h2;
parameter DDR_DDRC_CFG_RAS_CFG_RAS = 'h26;
parameter DDR_DDRC_CFG_RCD_CFG_RCD = 'hC;
parameter DDR_DDRC_CFG_RRD_CFG_RRD = 'h7;
parameter DDR_DDRC_CFG_RP_CFG_RP = 'hC;
parameter DDR_DDRC_CFG_RC_CFG_RC = 'h32;
parameter DDR_DDRC_CFG_FAW_CFG_FAW = 'h1B;
parameter DDR_DDRC_CFG_RFC_CFG_RFC = 'h76;
parameter DDR_DDRC_CFG_RTP_CFG_RTP = 'h8;
parameter DDR_DDRC_CFG_WR_CFG_WR = 'h10;
parameter DDR_DDRC_CFG_REF_PER_CFG_REF_PER = 'h207C;
parameter DDR_DDRC_CFG_STARTUP_DELAY_CFG_STARTUP_DELAY = 'hC8;
parameter DDR_DDRC_CFG_ZQ_CAL_PER_CFG_ZQ_CAL_PER = 'h3F40;
parameter DDR_DDRC_CFG_WTR_CFG_WTR = 'h8;
parameter DDR_DDRC_CFG_MOD_CFG_MOD = 'h10;
parameter DDR_DDRC_CFG_XS_CFG_XS = 'h80;
parameter DDR_DDRC_CFG_XPR_CFG_XPR = 'h80;
parameter DDR_DDRC_CFG_MANUAL_ADDRESS_MAP_CFG_MANUAL_ADDRESS_MAP = 'h0;
parameter DDR_DDRC_CFG_LOOKAHEAD_PCH_CFG_LOOKAHEAD_PCH = 'h1;
parameter DDR_DDRC_CFG_LOOKAHEAD_ACT_CFG_LOOKAHEAD_ACT = 'h1;
parameter DDR_DDRC_CFG_AUTO_REF_EN_CFG_AUTO_REF_EN = 'h1;
parameter DDR_DDRC_PHY_PC_RANK_PHY_PC_RANK = 'h0;
parameter DDR_DDRC_PHY_RANKS_TO_TRAIN_PHY_RANKS_TO_TRAIN = 'h3;
parameter DDR_DDRC_CFG_RMW_EN_CFG_RMW_EN = 'h1;
parameter DDR_DDRC_CFG_ECC_CORRECTION_EN_CFG_ECC_CORRECTION_EN = 'h1;
parameter DDR_DDRC_CFG_ONLY_SRANK_CMDS_CFG_ONLY_SRANK_CMDS = 'h0;
parameter DDR_DDRC_INIT_RDIMM_COMPLETE_INIT_RDIMM_COMPLETE = 'h0;
parameter DDR_DDRC_CFG_DM_EN_CFG_DM_EN = 'h1;
parameter DDR_DDRC_CFG_AL_MODE_CFG_AL_MODE = 'h0;
parameter DDR_DDRC_CFG_BL_MODE_CFG_BL_MODE = 'h0;
parameter DDR_DDRC_CFG_RTT_WR_CFG_RTT_WR = 'h0;
parameter DDR_DDRC_CFG_SRT_CFG_SRT = 'h0;
parameter DDR_DDRC_CFG_ADDR_MIRROR_CFG_ADDR_MIRROR = 'h0;
parameter DDR_DDRC_CFG_ZQ_CAL_TYPE_CFG_ZQ_CAL_TYPE = 'h0;
parameter DDR_DDRC_CFG_REGDIMM_CFG_REGDIMM = 'h0;
parameter DDR_DDRC_CFG_PASR_CFG_PASR = 'h0;
parameter DDR_DDRC_CFG_BT_CFG_BT = 'h0;
parameter DDR_DDRC_CFG_DS_CFG_DS = 'h0;
parameter DDR_DDRC_CFG_RTT_CFG_RTT = 'h1;
parameter DDR_DDRC_CFG_BANKADDR_MAP_1_CFG_BANKADDR_MAP_1 = 'h0;
parameter DDR_DDRC_CFG_NIBBLE_DEVICES_CFG_NIBBLE_DEVICES = 'h0;
parameter DDR_DDRC_CTRLR_SOFT_RESET_N_CTRLR_SOFT_RESET_N = 'h0;
parameter DDR_DDRC_CFG_READ_TO_WRITE_CFG_READ_TO_WRITE = 'h2;
parameter DDR_DDRC_CFG_WRITE_TO_WRITE_CFG_WRITE_TO_WRITE = 'h3;
parameter DDR_DDRC_CFG_READ_TO_READ_CFG_READ_TO_READ = 'h3;
parameter DDR_DDRC_CFG_WRITE_TO_READ_CFG_WRITE_TO_READ = 'h8;
parameter DDR_DDRC_CFG_READ_TO_WRITE_ODT_CFG_READ_TO_WRITE_ODT = 'h2;
parameter DDR_DDRC_CFG_WRITE_TO_WRITE_ODT_CFG_WRITE_TO_WRITE_ODT = 'h3;
parameter DDR_DDRC_CFG_READ_TO_READ_ODT_CFG_READ_TO_READ_ODT = 'h3;
parameter DDR_DDRC_CFG_WRITE_TO_READ_ODT_CFG_WRITE_TO_READ_ODT = 'h2;
parameter DDR_DDRC_CFG_MIN_READ_IDLE_CFG_MIN_READ_IDLE = 'h0;
parameter DDR_DDRC_CFG_QOFF_CFG_QOFF = 'h0;
parameter DDR_DDRC_CFG_DLL_DISABLE_CFG_DLL_DISABLE = 'h0;
parameter DDR_DDRC_CFG_ODT_RD_MAP_CS2_CFG_ODT_RD_MAP_CS2 = 'h8;
parameter DDR_DDRC_CFG_ODT_RD_MAP_CS3_CFG_ODT_RD_MAP_CS3 = 'h4;
parameter DDR_DDRC_CFG_ODT_RD_MAP_CS4_CFG_ODT_RD_MAP_CS4 = 'h20;
parameter DDR_DDRC_CFG_ODT_RD_MAP_CS5_CFG_ODT_RD_MAP_CS5 = 'h10;
parameter DDR_DDRC_CFG_ODT_RD_MAP_CS6_CFG_ODT_RD_MAP_CS6 = 'h80;
parameter DDR_DDRC_CFG_ODT_RD_MAP_CS7_CFG_ODT_RD_MAP_CS7 = 'h40;
parameter DDR_DDRC_CFG_ODT_WR_MAP_CS2_CFG_ODT_WR_MAP_CS2 = 'h4;
parameter DDR_DDRC_CFG_ODT_WR_MAP_CS3_CFG_ODT_WR_MAP_CS3 = 'h8;
parameter DDR_DDRC_CFG_ODT_WR_MAP_CS4_CFG_ODT_WR_MAP_CS4 = 'h10;
parameter DDR_DDRC_CFG_ODT_WR_MAP_CS5_CFG_ODT_WR_MAP_CS5 = 'h20;
parameter DDR_DDRC_CFG_ODT_WR_MAP_CS6_CFG_ODT_WR_MAP_CS6 = 'h40;
parameter DDR_DDRC_CFG_ODT_WR_MAP_CS7_CFG_ODT_WR_MAP_CS7 = 'h80;
parameter DDR_DDRC_CFG_ODT_RD_TURN_ON_CFG_ODT_RD_TURN_ON = 'h0;
parameter DDR_DDRC_CFG_ODT_WR_TURN_ON_CFG_ODT_WR_TURN_ON = 'h0;
parameter DDR_DDRC_CFG_ODT_RD_TURN_OFF_CFG_ODT_RD_TURN_OFF = 'h0;
parameter DDR_DDRC_CFG_ODT_WR_TURN_OFF_CFG_ODT_WR_TURN_OFF = 'h0;
parameter DDR_DDRC_CFG_EMR3_CFG_EMR3 = 'h0;
parameter DDR_DDRC_CFG_TWO_T_CFG_TWO_T = 'h0;
parameter DDR_DDRC_CFG_TWO_T_SEL_CYCLE_CFG_TWO_T_SEL_CYCLE = 'h0;
parameter DDR_DDRC_CFG_TDQS_CFG_TDQS = 'h0;
parameter DDR_DDRC_CFG_AUTO_SR_CFG_AUTO_SR = 'h0;
parameter DDR_DDRC_CFG_AUTO_ZQ_CAL_EN_CFG_AUTO_ZQ_CAL_EN = 'h1;
parameter DDR_DDRC_CFG_MEMORY_TYPE_CFG_MEMORY_TYPE = 'h8;
parameter DDR_DDRC_CFG_QUAD_RANK_CFG_QUAD_RANK = 'h0;
parameter DDR_DDRC_CFG_EARLY_RANK_TO_WR_START_CFG_EARLY_RANK_TO_WR_START = 'h0;
parameter DDR_DDRC_CFG_EARLY_RANK_TO_RD_START_CFG_EARLY_RANK_TO_RD_START = 'h0;
parameter DDR_DDRC_CFG_CAL_READ_PERIOD_CFG_CAL_READ_PERIOD = 'h0;
parameter DDR_DDRC_CFG_NUM_CAL_READS_CFG_NUM_CAL_READS = 'h0;
parameter DDR_DDRC_CFG_CTRLR_INIT_DISABLE_CFG_CTRLR_INIT_DISABLE = 'h0;
parameter DDR_DDRC_CFG_RDIMM_LAT_CFG_RDIMM_LAT = 'h0;
parameter DDR_DDRC_CFG_CTRLUPD_TRIG_CFG_CTRLUPD_TRIG = 'h1;
parameter DDR_DDRC_CFG_CTRLUPD_START_DELAY_CFG_CTRLUPD_START_DELAY = 'h16;
parameter DDR_DDRC_CFG_DFI_T_CTRLUPD_MAX_CFG_DFI_T_CTRLUPD_MAX = 'hC8;
parameter DDR_DDRC_CFG_DFI_T_RDDATA_EN_CFG_DFI_T_RDDATA_EN = 'h11;
parameter DDR_DDRC_CFG_DFI_T_PHY_WRLAT_CFG_DFI_T_PHY_WRLAT = 'h5;
parameter DDR_DDRC_PHY_DFI_INIT_START_PHY_DFI_INIT_START = 'h0;
parameter DDR_DDRC_PHY_RESET_CONTROL_PHY_RESET_CONTROL = 'h800D;
parameter DDR_DDRC_PHY_GATE_TRAIN_DELAY_PHY_GATE_TRAIN_DELAY = 'h1E;
parameter DDR_DDRC_PHY_EYE_TRAIN_DELAY_PHY_EYE_TRAIN_DELAY = 'h28;
parameter DDR_DDRC_PHY_TRAIN_STEP_ENABLE_PHY_TRAIN_STEP_ENABLE = 'h18;
parameter DDR_DDRC_PHY_INDPNDT_TRAINING_PHY_INDPNDT_TRAINING = 'h0;
parameter DDR_DDRC_CFG_DQ_WIDTH_CFG_DQ_WIDTH = 'h0;
parameter DDR_DDRC_CFG_CA_PARITY_ERR_STATUS_CFG_CA_PARITY_ERR_STATUS = 'h0;
parameter DDR_DDRC_CFG_PARITY_RDIMM_DELAY_CFG_PARITY_RDIMM_DELAY = 'h1;
parameter DDR_DDRC_CFG_DFI_T_PHY_RDLAT_CFG_DFI_T_PHY_RDLAT = 'h6;
parameter DDR_DDRC_CFG_DATA_MASK_CFG_DATA_MASK = 'h4;
parameter DDR_MODEL_DATA_LANES_USED_DATA_LANES = 'h4;
parameter DDR_DDRC_CFG_CCD_S_CFG_CCD_S = 'h5;
parameter DDR_DDRC_CFG_CCD_L_CFG_CCD_L = 'h6;
parameter DDR_DDRC_CFG_RRD_S_CFG_RRD_S = 'h4;
parameter DDR_DDRC_CFG_RRD_L_CFG_RRD_L = 'h3;
parameter DDR_DDRC_CFG_WTR_S_CFG_WTR_S = 'h3;
parameter DDR_DDRC_CFG_WTR_L_CFG_WTR_L = 'h3;
parameter DDR_DDRC_CFG_WTR_S_CRC_DM_CFG_WTR_S_CRC_DM = 'h3;
parameter DDR_DDRC_CFG_WTR_L_CRC_DM_CFG_WTR_L_CRC_DM = 'h3;
parameter DDR_DDRC_CFG_WR_CRC_DM_CFG_WR_CRC_DM = 'h6;
parameter DDR_DDRC_CFG_VREFDQ_TRN_VALUE_CFG_VREFDQ_TRN_VALUE = 'h0;
parameter DDR_DDRC_CFG_RFC1_CFG_RFC1 = 'h36;
parameter DDR_DDRC_CFG_RFC2_CFG_RFC2 = 'h36;
parameter DDR_DDRC_CFG_RFC4_CFG_RFC4 = 'h36;
parameter DDR_DDRC_CFG_FINE_GRAN_REF_MODE_CFG_FINE_GRAN_REF_MODE = 'h0;
parameter DDR_DDRC_CFG_RD_PREAMBLE_CFG_RD_PREAMBLE = 'h0;
parameter DDR_DDRC_CFG_SR_ABORT_CFG_SR_ABORT = 'h0;
parameter DDR_DDRC_CFG_INT_VREF_MON_CFG_INT_VREF_MON = 'h0;
parameter DDR_DDRC_CFG_TEMP_CTRL_REF_MODE_CFG_TEMP_CTRL_REF_MODE = 'h0;
parameter DDR_DDRC_CFG_TEMP_CTRL_REF_RANGE_CFG_TEMP_CTRL_REF_RANGE = 'h0;
parameter DDR_DDRC_CFG_RTT_PARK_CFG_RTT_PARK = 'h0;
parameter DDR_DDRC_CFG_ODT_INBUF_4_PD_CFG_ODT_INBUF_4_PD = 'h0;
parameter DDR_DDRC_CFG_CA_PARITY_LATENCY_CFG_CA_PARITY_LATENCY = 'h0;
parameter DDR_DDRC_CFG_VREFDQ_TRN_ENABLE_CFG_VREFDQ_TRN_ENABLE = 'h0;
parameter DDR_DDRC_CFG_VREFDQ_TRN_RANGE_CFG_VREFDQ_TRN_RANGE = 'h0;
parameter DDR_DDRC_CFG_LP_ASR_CFG_LP_ASR = 'h0;
parameter DDR_DDRC_CFG_WR_PREAMBLE_CFG_WR_PREAMBLE = 'h0;
parameter DDR_DDRC_CFG_RFC_DLR1_CFG_RFC_DLR1 = 'h48;
parameter DDR_DDRC_CFG_RFC_DLR2_CFG_RFC_DLR2 = 'h2C;
parameter DDR_DDRC_CFG_RFC_DLR4_CFG_RFC_DLR4 = 'h20;
parameter DDR_DDRC_CFG_RRD_DLR_CFG_RRD_DLR = 'h4;
parameter DDR_DDRC_CFG_FAW_DLR_CFG_FAW_DLR = 'h10;
parameter DDR_DDRC_CFG_BG_INTERLEAVE_CFG_BG_INTERLEAVE = 'h1;
parameter DDR_DDRC_CFG_MRR_CFG_MRR = 'h2;
parameter DDR_DDRC_CFG_MRW_CFG_MRW = 'h10;
parameter DDR_DDRC_CFG_XP_CFG_XP = 'h3;
parameter DDR_DDRC_CFG_XSR_CFG_XSR = 'h24;
parameter DDR_DDRC_CFG_INIT_DURATION_CFG_INIT_DURATION = 'h29B0;
parameter DDR_DDRC_CFG_ZQ_CAL_R_DURATION_CFG_ZQ_CAL_R_DURATION = 'hB;
parameter DDR_DDRC_CFG_ODT_POWERDOWN_CFG_ODT_POWERDOWN = 'h0;
parameter DDR_DDRC_CFG_WL_CFG_WL = 'h9;
parameter DDR_DDRC_CFG_RL_CFG_RL = 'hC;
parameter DDR_DDRC_CFG_BL_CFG_BL = 'h0;
parameter DDR_OPTIONS_TIP_CFG_PARAMS_ADDCMD_OFFSET = 'h0;
parameter DDR_DDRC_CFG_ZQLATCH_DURATION_CFG_ZQLATCH_DURATION = 'h30;
parameter DDR_DDRC_CFG_ZQ_CAL_DURATION_CFG_ZQ_CAL_DURATION = 'h640;
parameter DDR_DDRC_CFG_MRRI_CFG_MRRI = 'h0;
parameter DDR_DDRC_CFG_WR_POSTAMBLE_CFG_WR_POSTAMBLE = 'h0;
parameter DDR_DDRC_CFG_SOC_ODT_CFG_SOC_ODT = 'h0;
parameter DDR_DDRC_CFG_ODTE_CK_CFG_ODTE_CK = 'h0;
parameter DDR_DDRC_CFG_ODTE_CS_CFG_ODTE_CS = 'h0;
parameter DDR_DDRC_CFG_ODTD_CA_CFG_ODTD_CA = 'h0;
parameter DDR_DDRC_CFG_RD_PREAMB_TOGGLE_CFG_RD_PREAMB_TOGGLE = 'h0;
parameter DDR_DDRC_CFG_RD_POSTAMBLE_CFG_RD_POSTAMBLE = 'h0;
parameter DDR_DDRC_CFG_PU_CAL_CFG_PU_CAL = 'h0;
parameter DDR_DDRC_CFG_DQ_ODT_CFG_DQ_ODT = 'h0;
parameter DDR_DDRC_CFG_CA_ODT_CFG_CA_ODT = 'h0;
parameter DDR_DDRC_CFG_MRD_CFG_MRD = 'h10;
parameter DDR_DDRC_CFG_LPDDR4_FSP_OP_CFG_LPDDR4_FSP_OP = 'h0;
parameter CLK_MSS_SYS_CLOCK_CONFIG_CR_DIVIDER_CPU = 'h0;
parameter CLK_MSS_SYS_CLOCK_CONFIG_CR_DIVIDER_AXI = 'h1;
parameter CLK_MSS_SYS_CLOCK_CONFIG_CR_DIVIDER_APB_AHB = 'h2;
parameter CLK_MSS_CFM_PLL_CKMUX_PLL1_RFCLK0_SEL = 'h1;
parameter CLK_MSS_CFM_PLL_CKMUX_PLL1_RFCLK1_SEL = 'h1;
parameter CLK_MSS_CFM_PLL_CKMUX_PLL0_RFCLK0_SEL = 'h1;
parameter CLK_MSS_CFM_PLL_CKMUX_PLL0_RFCLK1_SEL = 'h1;
parameter CLK_MSS_CFM_PLL_CKMUX_CLK_IN_MAC_TSU_SEL = 'h1;
parameter SGMII_CLK_CNTL_REG_CLKMUX_PLL0_RFCLK0_SEL = 'h1;
parameter SGMII_CLK_CNTL_REG_CLKMUX_PLL0_RFCLK1_SEL = 'h1;
parameter CLK_MSS_CFM_MSSCLKMUX_MSSCLK_MUX_SEL = 'h3;
parameter CLK_MSS_CFM_MSSCLKMUX_CLK_STANDBY_SEL = 'h0;
parameter CLK_MSS_CFM_BCLKMUX_BCLK0_SEL = 'h8;
parameter CLK_MSS_CFM_BCLKMUX_BCLK1_SEL = 'h10;
parameter CLK_MSS_CFM_BCLKMUX_BCLK2_SEL = 'h0;
parameter CLK_MSS_CFM_BCLKMUX_BCLK3_SEL = 'h0;
parameter CLK_MSS_CFM_BCLKMUX_BCLK4_SEL = 'h0;
parameter CLK_MSS_CFM_BCLKMUX_BCLK5_SEL = 'h0;
parameter CLK_MSS_PLL_PLL_CTRL_REG_RFCLK_SEL = 'h0;
parameter CLK_SGMII_PLL_PLL_CTRL_REG_RFCLK_SEL = 'h0;
parameter CLK_DDR_PLL_PLL_CTRL_REG_RFCLK_SEL = 'h0;
parameter DDR_MODEL_DDRPHY_MODE_DDRMODE = 'h7;
parameter DDR_MODEL_DDRPHY_MODE_POWER_DOWN = 'h1;
parameter DDR_MODEL_DDRPHY_MODE_CRC = 'h0;
parameter DDR_MODEL_DDRPHY_MODE_ECC = 'h1;
parameter DDR_MODEL_DDRPHY_MODE_BUS_WIDTH = 'h1;
parameter DDR_MODEL_DDRPHY_MODE_DMI_DBI = 'h1;
parameter DDR_MODEL_DDRPHY_MODE_RANK = 'h1;
parameter DDR_MODEL_DDRPHY_MODE_DQ_DRIVE = 'h0;
parameter DDR_MODEL_DDRPHY_MODE_DQS_DRIVE = 'h0;
parameter DDR_MODEL_DDRPHY_MODE_ADD_CMD_DRIVE = 'h0;
parameter DDR_MODEL_DDRPHY_MODE_CLOCK_OUT_DRIVE = 'h0;
parameter DDR_IOBANK_RPC_ODT_DQ_RPC_ODT_DQ = 'h4;
parameter DDR_IOBANK_RPC_ODT_DQS_RPC_ODT_DQS = 'h4;
parameter DDR_IOBANK_DPC_BITS_DPC_VRGEN_V = 'h1E;
parameter DDR_IOBANK_DPC_BITS_DPC_VRGEN_H = 'h3C;
parameter DDR_IOBANK_DPC_BITS_DPC_VRGEN_EN_V = 'h1;
parameter DDR_IOBANK_DPC_BITS_DPC_VRGEN_EN_H = 'h1;
parameter DDR_IOBANK_DPC_BITS_DPC_MOVE_EN_V = 'h0;
parameter DDR_IOBANK_DPC_BITS_DPC_MOVE_EN_H = 'h0;
parameter DDR_IOBANK_DPC_BITS_DPC_VS = 'h5;
parameter DDR_IOBANK_RPC_ODT_STATIC_DQ_RPC_ODT_STATIC_DQ = 'h7;
parameter DDR_IOBANK_RPC_ODT_STATIC_DQS_RPC_ODT_STATIC_DQS = 'h7;
parameter DDR_IOBANK_RPC_ODT_STATIC_ADDCMD_RPC_ODT_STATIC_ADDCMD = 'h7;
parameter DDR_IOBANK_RPC_ODT_STATIC_CLKP_RPC_ODT_STATIC_CLKP = 'h7;
parameter DDR_IOBANK_RPC_ODT_STATIC_CLKN_RPC_ODT_STATIC_CLKN = 'h7;
parameter DDR_IOBANK_RPC_IBUFMD_ADDCMD_RPC_IBUFMD_ADDCMD = 'h3;
parameter DDR_IOBANK_RPC_IBUFMD_CLK_RPC_IBUFMD_CLK = 'h4;
parameter DDR_IOBANK_RPC_IBUFMD_DQ_RPC_IBUFMD_DQ = 'h3;
parameter DDR_IOBANK_RPC_IBUFMD_DQS_RPC_IBUFMD_DQS = 'h4;
parameter DDR_IOBANK_RPC_SPARE0_DQ_RPC_SPARE0_DQ = 'h0;
parameter SGMII_SPARE_CNTL_REG_SPARE = 'h0;
parameter TRACE_CR_ULTRASOC_FABRIC = 'h0;
parameter MSS_IO_LOCKDOWN_CR_MSSIO_B2_LOCKDN_EN = 'h0;
parameter MSS_IO_LOCKDOWN_CR_MSSIO_B4_LOCKDN_EN = 'h0;
parameter MSS_IO_LOCKDOWN_CR_SGMII_IO_LOCKDN_EN = 'h0;
parameter MSS_IO_LOCKDOWN_CR_DDR_IO_LOCKDN_EN = 'h0;
parameter DLL0_CTRL0_PHASE_P = 'h0;
parameter DLL0_CTRL0_PHASE_S = 'h0;
parameter DLL0_CTRL0_SEL_P = 'h0;
parameter DLL0_CTRL0_SEL_S = 'h0;
parameter DLL0_CTRL0_REF_SEL = 'h0;
parameter DLL0_CTRL0_FB_SEL = 'h0;
parameter DLL0_CTRL0_DIV_SEL = 'h0;
parameter DLL0_CTRL0_ALU_UPD = 'h0;
parameter DLL0_CTRL0_LOCK_FRC = 'h0;
parameter DLL0_CTRL0_LOCK_FLT = 'h0;
parameter DLL0_CTRL0_LOCK_HIGH = 'h0;
parameter DLL0_CTRL0_LOCK_LOW = 'h0;
parameter DLL0_CTRL1_SET_ALU = 'h0;
parameter DLL0_CTRL1_ADJ_DEL4 = 'h0;
parameter DLL0_CTRL1_TEST_S = 'h0;
parameter DLL0_CTRL1_TEST_RING = 'h0;
parameter DLL0_CTRL1_INIT_CODE = 'h0;
parameter DLL0_CTRL1_RELOCK_FAST = 'h0;
parameter DLL0_STAT0_RESET = 'h0;
parameter DLL0_STAT0_BYPASS = 'h0;
parameter DLL0_STAT0_PHASE_MOVE_CLK = 'h0;
parameter DLL1_CTRL0_PHASE_P = 'h0;
parameter DLL1_CTRL0_PHASE_S = 'h0;
parameter DLL1_CTRL0_SEL_P = 'h0;
parameter DLL1_CTRL0_SEL_S = 'h0;
parameter DLL1_CTRL0_REF_SEL = 'h0;
parameter DLL1_CTRL0_FB_SEL = 'h0;
parameter DLL1_CTRL0_DIV_SEL = 'h0;
parameter DLL1_CTRL0_ALU_UPD = 'h0;
parameter DLL1_CTRL0_LOCK_FRC = 'h0;
parameter DLL1_CTRL0_LOCK_FLT = 'h0;
parameter DLL1_CTRL0_LOCK_HIGH = 'h0;
parameter DLL1_CTRL0_LOCK_LOW = 'h0;
parameter DLL1_CTRL1_SET_ALU = 'h0;
parameter DLL1_CTRL1_ADJ_DEL4 = 'h0;
parameter DLL1_CTRL1_TEST_S = 'h0;
parameter DLL1_CTRL1_TEST_RING = 'h0;
parameter DLL1_CTRL1_INIT_CODE = 'h0;
parameter DLL1_CTRL1_RELOCK_FAST = 'h0;
parameter DLL1_STAT0_RESET = 'h0;
parameter DLL1_STAT0_BYPASS = 'h0;
parameter DLL1_STAT0_PHASE_MOVE_CLK = 'h0;
parameter DLL2_CTRL0_PHASE_P = 'h0;
parameter DLL2_CTRL0_PHASE_S = 'h0;
parameter DLL2_CTRL0_SEL_P = 'h0;
parameter DLL2_CTRL0_SEL_S = 'h0;
parameter DLL2_CTRL0_REF_SEL = 'h0;
parameter DLL2_CTRL0_FB_SEL = 'h0;
parameter DLL2_CTRL0_DIV_SEL = 'h0;
parameter DLL2_CTRL0_ALU_UPD = 'h0;
parameter DLL2_CTRL0_LOCK_FRC = 'h0;
parameter DLL2_CTRL0_LOCK_FLT = 'h0;
parameter DLL2_CTRL0_LOCK_HIGH = 'h0;
parameter DLL2_CTRL0_LOCK_LOW = 'h0;
parameter DLL2_CTRL1_SET_ALU = 'h0;
parameter DLL2_CTRL1_ADJ_DEL4 = 'h0;
parameter DLL2_CTRL1_TEST_S = 'h0;
parameter DLL2_CTRL1_TEST_RING = 'h0;
parameter DLL2_CTRL1_INIT_CODE = 'h0;
parameter DLL2_CTRL1_RELOCK_FAST = 'h0;
parameter DLL2_STAT0_RESET = 'h0;
parameter DLL2_STAT0_BYPASS = 'h0;
parameter DLL2_STAT0_PHASE_MOVE_CLK = 'h0;
parameter DLL3_CTRL0_PHASE_P = 'h0;
parameter DLL3_CTRL0_PHASE_S = 'h0;
parameter DLL3_CTRL0_SEL_P = 'h0;
parameter DLL3_CTRL0_SEL_S = 'h0;
parameter DLL3_CTRL0_REF_SEL = 'h0;
parameter DLL3_CTRL0_FB_SEL = 'h0;
parameter DLL3_CTRL0_DIV_SEL = 'h0;
parameter DLL3_CTRL0_ALU_UPD = 'h0;
parameter DLL3_CTRL0_LOCK_FRC = 'h0;
parameter DLL3_CTRL0_LOCK_FLT = 'h0;
parameter DLL3_CTRL0_LOCK_HIGH = 'h0;
parameter DLL3_CTRL0_LOCK_LOW = 'h0;
parameter DLL3_CTRL1_SET_ALU = 'h0;
parameter DLL3_CTRL1_ADJ_DEL4 = 'h0;
parameter DLL3_CTRL1_TEST_S = 'h0;
parameter DLL3_CTRL1_TEST_RING = 'h0;
parameter DLL3_CTRL1_INIT_CODE = 'h0;
parameter DLL3_CTRL1_RELOCK_FAST = 'h0;
parameter DLL3_STAT0_RESET = 'h0;
parameter DLL3_STAT0_BYPASS = 'h0;
parameter DLL3_STAT0_PHASE_MOVE_CLK = 'h0;
parameter CRYPTO_SOFT_RESET_PERIPH = 'h0;
parameter CRYPTO_DLL_CTRL0_PHASE_P = 'h0;
parameter CRYPTO_DLL_CTRL0_PHASE_S = 'h0;
parameter CRYPTO_DLL_CTRL0_SEL_P = 'h0;
parameter CRYPTO_DLL_CTRL0_SEL_S = 'h0;
parameter CRYPTO_DLL_CTRL0_REF_SEL = 'h0;
parameter CRYPTO_DLL_CTRL0_FB_SEL = 'h0;
parameter CRYPTO_DLL_CTRL0_DIV_SEL = 'h0;
parameter CRYPTO_DLL_CTRL0_ALU_UPD = 'h0;
parameter CRYPTO_DLL_CTRL0_LOCK_FRC = 'h0;
parameter CRYPTO_DLL_CTRL0_LOCK_FLT = 'h0;
parameter CRYPTO_DLL_CTRL0_LOCK_HIGH = 'h0;
parameter CRYPTO_DLL_CTRL0_LOCK_LOW = 'h0;
parameter CRYPTO_DLL_CTRL1_SET_ALU = 'h0;
parameter CRYPTO_DLL_CTRL1_ADJ_DEL4 = 'h0;
parameter CRYPTO_DLL_CTRL1_TEST_S = 'h0;
parameter CRYPTO_DLL_CTRL1_TEST_RING = 'h0;
parameter CRYPTO_DLL_CTRL1_INIT_CODE = 'h0;
parameter CRYPTO_DLL_CTRL1_RELOCK_FAST = 'h0;
parameter CRYPTO_DLL_STAT0_RESET = 'h0;
parameter CRYPTO_DLL_STAT0_BYPASS = 'h0;
parameter CRYPTO_DLL_STAT0_PHASE_MOVE_CLK = 'h0;
parameter CRYPTO_CONTROL_USER_SCB_CONTROL = 'h0;
parameter CRYPTO_CONTROL_USER_RESET = 'h0;
parameter CRYPTO_CONTROL_USER_CLOCK_ENABLE = 'h0;
parameter CRYPTO_CONTROL_USER_CLOCK_SELECT = 'h0;
parameter CRYPTO_CONTROL_USER_RAMS_ON = 'h0;
parameter CRYPTO_CONTROL_USER_DLL_ON = 'h0;
parameter CRYPTO_CONTROL_USER_RING_OSC_ON = 'h0;
parameter CRYPTO_CONTROL_USER_PURGE = 'h0;
parameter CRYPTO_CONTROL_USER_GO = 'h0;
parameter CRYPTO_INTERRUPT_ENABLE_COMPLETE = 'h0;
parameter CRYPTO_INTERRUPT_ENABLE_ALARM = 'h0;
parameter CRYPTO_INTERRUPT_ENABLE_BUSERROR = 'h0;
parameter CRYPTO_MARGIN_RAM = 'h0;
parameter CRYPTO_MARGIN_ROM = 'h0;

endmodule
